//Constant array to load the A matrix
localparam integer A_size = 11;
localparam integer A[0:10] = '{32'h40a00000, 32'h40000000, 32'h3f800000, 32'h40800000, 32'hc0400000, 32'hc0a00000, 32'hc0000000, 32'hc0800000, 32'hbf800000, 32'h40c00000, 32'h40400000};
localparam integer A_BRAMInd[0:10] = '{0, 1, 2, 3, 0, 1, 0, 1, 2, 3, 2};
localparam integer A_BRAMAddr[0:10] = '{0, 0, 0, 0, 1, 1, 2, 2, 2, 2, 3};

//Constant array to load the instruction BRAM
localparam integer total_instructions = 54;
localparam integer sub_instructions = 3;
localparam integer Inst[0:53][0:2] = '{{32'h0, 32'h0, 32'h0},{32'h34000, 32'h80000, 32'h0},{32'h44c00, 32'h20000000, 32'h1},{32'h0, 32'h40000000, 32'h0},{32'h2a000, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h1},{32'h44700080, 32'h40000, 32'h0},{32'h4a700010, 32'h80, 32'h0},{32'haf00000, 32'h100200, 32'h0},{32'h6600400, 32'h60080000, 32'h0},{32'h7300000, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h80000000, 32'h0},{32'h20000, 32'h180, 32'h0},{32'h0, 32'h1c0000, 32'h0},{32'h70000000, 32'he0000000, 32'h0},{32'h0, 32'h280, 32'h0},{32'h30000000, 32'h0, 32'h0},{32'h20000000, 32'h100, 32'h0},{32'h58000, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h60000000, 32'h300, 32'h0},{32'ha600400, 32'ha0000000, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h30000002, 32'h0, 32'h0},{32'h20000000, 32'hc0180000, 32'h0},{32'h5580000, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h380, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h1c0000, 32'h0},{32'h0, 32'h0, 32'h0},{32'h1, 32'h0, 32'h0}};

