//Constant array to load the A matrix
localparam integer A_size = 10;
localparam integer A[0:9] = '{32'h41000000, 32'h3f800000, 32'h40e00000, 32'h40a00000, 32'h40000000, 32'hc0000000, 32'h3f800000, 32'h40000000, 32'hc0400000, 32'h41100000};
localparam integer A_BRAMInd[0:9] = '{0, 1, 0, 1, 1, 0, 1, 0, 1, 0};
localparam integer A_BRAMAddr[0:9] = '{0, 0, 1, 1, 2, 3, 3, 5, 5, 6};

//Constant array to load the instruction BRAM
localparam integer total_instructions = 161;
localparam integer sub_instructions = 2;
localparam integer Inst[0:160][0:1] = '{{32'h60000000, 32'h0},{32'h20045400, 32'hf00040},{32'h4a000, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h200000},{32'h4700010, 32'he00010},{32'h4700010, 32'h600050},{32'h5700000, 32'hc0a040},{32'h7100000, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h20},{32'h8000, 32'h0},{32'h0, 32'h90},{32'h0, 32'h900000},{32'h0, 32'hd00000},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'ha000a0},{32'h4600400, 32'h500000},{32'h0, 32'h804060},{32'h8d00000, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'hb0},{32'h0, 32'h80},{32'h40000, 32'h900000},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h10, 32'h90},{32'h80000000, 32'hc000a0},{32'h9500000, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'h0},{32'h0, 32'hd00000},{32'h0, 32'h0},{32'h1, 32'h0}};

