//Constant array to load the A matrix
localparam integer A_size = 665;
localparam integer A[0:664] = '{32'h3e088c61, 32'hbd8888b5, 32'hb76ae18b, 32'hbd8888b5, 32'h3e088c61, 32'hbd8888b5, 32'hb76ae18b, 32'hbd8888b5, 32'h3e088ace, 32'hbd8888b5, 32'hbd8888b5, 32'hb70637bd, 32'h4170021b, 32'hb9fa9c13, 32'hb58637bd, 32'hb796feb5, 32'hb796feb5, 32'hb9fb224b, 32'h3b272eae, 32'hb8b88ca4, 32'hba828c37, 32'hba81a155, 32'hbd8888b5, 32'hbd8888b5, 32'h360637bd, 32'h390b75ea, 32'h3eaad2fe, 32'hb9712c28, 32'hbe4ccccd, 32'hb95f58c1, 32'hb76ae18b, 32'hb78637bd, 32'hbab02928, 32'h39ad8a11, 32'h3c51dcd7, 32'hbc441dd2, 32'h3955e8d5, 32'h3e08900c, 32'hbd8888b5, 32'hb7f34507, 32'hbd8888b5, 32'h3e088bdb, 32'hbd8888b5, 32'hbd8888b5, 32'hb75a1a93, 32'h40f00560, 32'hba19e0e7, 32'hb58637bd, 32'hb816feb5, 32'hb80a697b, 32'hba1aaa3b, 32'h3b81450f, 32'hba2d46f6, 32'hbad6909b, 32'hba8a8b09, 32'hbd8888b5, 32'hbd8888b5, 32'h368637bd, 32'h3948472c, 32'h3eaae4d2, 32'hb9d23d4f, 32'hbe4ccccd, 32'hb9798fa3, 32'hb7f34507, 32'hb81f6230, 32'hbb6874c9, 32'h3966afcd, 32'h3cd55821, 32'hbcc41dd2, 32'h3aa91538, 32'h3e088c61, 32'hb76ae18b, 32'hbd8888b5, 32'h3e088ace, 32'hbd8888b5, 32'hb716feb5, 32'h3cf3c2db, 32'hb87fda40, 32'hb58637bd, 32'hbcf2c301, 32'hb87fda40, 32'hb76ae18b, 32'hb8a5accd, 32'h3c69680e, 32'h3851b717, 32'hb78e9b39, 32'hbb113a50, 32'hbd8888b5, 32'hbd8888b5, 32'h36c9539c, 32'hb76ae18b, 32'h3eaaad1d, 32'h358637bd, 32'hb749539c, 32'hbcf2c301, 32'hb796feb5, 32'h3f5cedc4, 32'hb796feb5, 32'hbf555550, 32'h3d13165d, 32'hbcc41dd2, 32'hbc441dd2, 32'h3e08900c, 32'hbd8888b5, 32'hbd8888b5, 32'hb7f34507, 32'h3f800000, 32'hbd8888b5, 32'h3e088bdb, 32'hbd8888b5, 32'hb75a1a93, 32'hbd8888b5, 32'hbe4ccccd, 32'hbd8888b5, 32'h3eaaaf14, 32'hb6a7c5ac, 32'hb80a697b, 32'h36a7c5ac, 32'hb7f34507, 32'hbcc41dd2, 32'h358637bd, 32'h3cc4d445, 32'hb58637bd, 32'hb80e9b39, 32'hb7c9539c, 32'hb80637bd, 32'hb79f6230, 32'h3b8c2614, 32'hbb8b08dd, 32'h378e9b39, 32'hb80e9b39, 32'hbb8b08dd, 32'h3ed78983, 32'hb7e27e0f, 32'hbed55561, 32'hbcc41dd2, 32'hb75a1a93, 32'hb60637bd, 32'hb7e27e0f, 32'h3cc475e6, 32'hb716feb5, 32'hb851b717, 32'hbb0e25c8, 32'hb88e9b39, 32'hb7a7c5ac, 32'hbc441dd2, 32'h3c6a0ba2, 32'h3f800000, 32'h3e088c61, 32'hb76ae18b, 32'hbd8888b5, 32'hb76ae18b, 32'h3c449fd8, 32'hb78637bd, 32'h3e088a48, 32'hbd8888b5, 32'hb6c9539c, 32'h3bd6c2f0, 32'hb716feb5, 32'hb727c5ac, 32'hbbd6238e, 32'hbd8888b5, 32'hbd8888b5, 32'hb79f6230, 32'h3eaaad1d, 32'hb6c9539c, 32'hb727c5ac, 32'h3c449ba6, 32'hb76ae18b, 32'hbc441dd2, 32'hbf555550, 32'hb78637bd, 32'hbbd6238e, 32'hb76ae18b, 32'h3f57038e, 32'h40055554, 32'hbf555550, 32'h3f800000, 32'hbed55561, 32'hbf555550, 32'hbd8888b5, 32'h3e08900c, 32'hbd8888b5, 32'hb7f34507, 32'hbd8888b5, 32'h3e088d2a, 32'hbd8888b5, 32'hb796feb5, 32'hbe4ccccd, 32'hbd8888b5, 32'hbd8888b5, 32'h3eaaaf79, 32'hb7da1a93, 32'h377ba882, 32'hb7da1a93, 32'hbcc41dd2, 32'hb7f34507, 32'h38e27e0f, 32'h3ccfd8f1, 32'hb910b418, 32'hbaaf5fd4, 32'hb812ccf7, 32'hb6c9539c, 32'hb8e8c8ac, 32'h3c8f861a, 32'hb8e8c8ac, 32'hbc8da7f4, 32'hb796feb5, 32'hb910b418, 32'hbaa15981, 32'hb8dc3372, 32'h3cd0a244, 32'hb816feb5, 32'hbcc41dd2, 32'hbed55561, 32'hb816feb5, 32'hbc8da7f4, 32'hb816feb5, 32'h3ede392e, 32'h3cc41dd2, 32'hbc441dd2, 32'hbc441dd2, 32'h3e088c61, 32'hb76ae18b, 32'hbd8888b5, 32'hbc441dd2, 32'hb76ae18b, 32'h3c449fd8, 32'hb78637bd, 32'h3e088a48, 32'hb6eae18b, 32'hbd8888b5, 32'h3bd66f0d, 32'hb60637bd, 32'hb78637bd, 32'hbbd5cfab, 32'hb6eae18b, 32'h3c447a18, 32'hb60637bd, 32'hb76ae18b, 32'hbc441dd2, 32'hbd8888b5, 32'hbd8888b5, 32'hb79f6230, 32'h3eaaad1d, 32'hbf555550, 32'hb78637bd, 32'hbbd5cfab, 32'hb76ae18b, 32'h3f5702f7, 32'h3e088c61, 32'hb76ae18b, 32'hbd8888b5, 32'h3e088ace, 32'hbd8888b5, 32'hb716feb5, 32'h3cf02c4d, 32'hb896feb5, 32'hb60637bd, 32'hbceef805, 32'hb8991794, 32'hb76ae18b, 32'hb8dc3372, 32'h3c698138, 32'h385a1a93, 32'hb77ba882, 32'hbb101d19, 32'hbd8888b5, 32'hbd8888b5, 32'h36c9539c, 32'hb77ba882, 32'h3eaaad1d, 32'h3649539c, 32'hb749539c, 32'h3e088c61, 32'hb76ae18b, 32'hbd8888b5, 32'hb76ae18b, 32'h3c449fd8, 32'hb78637bd, 32'h3e088a48, 32'hbd8888b5, 32'hb6c9539c, 32'h3bd6ba8c, 32'hb727c5ac, 32'hb716feb5, 32'hbbd6238e, 32'hbd8888b5, 32'hbd8888b5, 32'hb79f6230, 32'h3eaaad1d, 32'hb6c9539c, 32'hb716feb5, 32'h3c449774, 32'hb76ae18b, 32'hbc441dd2, 32'hb78637bd, 32'hbbd6238e, 32'hb76ae18b, 32'h3f57038e, 32'hbf555550, 32'h3f800000, 32'h3e088c61, 32'hb76ae18b, 32'hbd8888b5, 32'hb76ae18b, 32'h3c449fd8, 32'hb78637bd, 32'h3bd6a9c5, 32'hb79f6230, 32'hbbd60a63, 32'h3e088a48, 32'hbd8888b5, 32'hb6eae18b, 32'hbd8888b5, 32'hb79f6230, 32'hbd8888b5, 32'h3eaaad1d, 32'hb6eae18b, 32'h3c4471b4, 32'hbc441dd2, 32'hb76ae18b, 32'hbc441dd2, 32'h3cc41dd2, 32'hbc441dd2, 32'hbf555550, 32'hb78637bd, 32'hbbd60a63, 32'hb76ae18b, 32'h3f57035c, 32'hbf555550, 32'h40055554, 32'hbf555550, 32'h3f800000, 32'hbed55561, 32'hbd8888b5, 32'h3e08900c, 32'hbd8888b5, 32'hb7f34507, 32'hbd8888b5, 32'h3e088d2a, 32'hbd8888b5, 32'hb796feb5, 32'hbe4ccccd, 32'hbd8888b5, 32'hbd8888b5, 32'h3eaaaf79, 32'hb7f34507, 32'h377ba882, 32'hb7c0f020, 32'hbcc41dd2, 32'hb7f34507, 32'h38e06530, 32'h3ccfce74, 32'hb910b418, 32'hbaae9681, 32'hb812ccf7, 32'hb6c9539c, 32'hb8e6afcd, 32'h3c8f1b26, 32'hb8e8c8ac, 32'hbc8d3cff, 32'hb796feb5, 32'hb910b418, 32'hbaa04d12, 32'hb8da1a93, 32'h3cd08f65, 32'hb816feb5, 32'hbcc41dd2, 32'hbed55561, 32'hb816feb5, 32'hbc8d3cff, 32'hb816feb5, 32'h3ede327f, 32'hbc441dd2, 32'hbcc41dd2, 32'h3f5e86b6, 32'hbf555550, 32'h3e088b54, 32'hbd8888b5, 32'hb7388ca4, 32'h3e088a48, 32'hbd8888b5, 32'hb6eae18b, 32'hbd8888b5, 32'hbd8888b5, 32'h3eaaac11, 32'hb727c5ac, 32'hb727c5ac, 32'h3b73eccc, 32'hbb734507, 32'h358637bd, 32'hb58637bd, 32'hbb734507, 32'h3f564ae0, 32'hb78e9b39, 32'hb78e9b39, 32'hbf555550, 32'hb6eae18b, 32'hb78e9b39, 32'h3c44827b, 32'hbc441dd2, 32'hbc441dd2, 32'hb7388ca4, 32'hb78e9b39, 32'hb58637bd, 32'h3c449774, 32'hbceef805, 32'hb796feb5, 32'hbf555550, 32'h3f5ccf5b, 32'hb796feb5, 32'hbc441dd2, 32'hb716feb5, 32'hb849539c, 32'hbb0dc11e, 32'hb890b418, 32'hb7b88ca4, 32'h3c69fadb, 32'hbc441dd2, 32'hbcc41dd2, 32'hbf555550, 32'h3f5e86b6, 32'hbc441dd2, 32'h3f5b763e, 32'hbf555550, 32'hbc441dd2, 32'h3e088c61, 32'hb76ae18b, 32'hbd8888b5, 32'h3e088ace, 32'hbd8888b5, 32'hb716feb5, 32'h3cf03afb, 32'hb88205ff, 32'hb58637bd, 32'hbcef3d3a, 32'hb8734507, 32'hb76ae18b, 32'hb8a17b0f, 32'h3c689a89, 32'h384d8559, 32'hb78e9b39, 32'hbb0e1501, 32'hbd8888b5, 32'hbd8888b5, 32'h36c9539c, 32'hb80a697b, 32'h3eaaacfb, 32'h358637bd, 32'h36eae18b, 32'hbcef3d3a, 32'hb796feb5, 32'h3f5cd196, 32'hb796feb5, 32'hbf555550, 32'h3d13165d, 32'hbc441dd2, 32'hbcc41dd2, 32'h3e088c61, 32'hbd8888b5, 32'hb76ae18b, 32'h3e088a48, 32'hbd8888b5, 32'hb6c9539c, 32'hbd8888b5, 32'hbd8888b5, 32'h3eaaacfb, 32'hb796feb5, 32'hb76ae18b, 32'h3c44a83b, 32'hb78e9b39, 32'hb60637bd, 32'hb75a1a93, 32'hb58637bd, 32'h3bd7a56e, 32'hbbd70e6f, 32'hb68637bd, 32'hb78e9b39, 32'hbbd70e6f, 32'h3f570564, 32'hb76ae18b, 32'hbf555550, 32'hbc441dd2, 32'hb6c9539c, 32'hb6a7c5ac, 32'hb76ae18b, 32'h3c4486ad, 32'hbd8888b5, 32'h3e08900c, 32'hbd8888b5, 32'hb7f34507, 32'hbd8888b5, 32'h3e088d2a, 32'hbd8888b5, 32'hb796feb5, 32'hbe4ccccd, 32'hbd8888b5, 32'hbd8888b5, 32'h3eaaaf79, 32'hb7da1a93, 32'h377ba882, 32'hb7da1a93, 32'hbcc41dd2, 32'hb7f34507, 32'h38dc3372, 32'h3ccfe154, 32'hb90d8ec9, 32'hbaafe60c, 32'hb816feb5, 32'hb68637bd, 32'hb8e8c8ac, 32'h3c90752e, 32'hb8e8c8ac, 32'hbc8e9d52, 32'hbcc41dd2, 32'hb796feb5, 32'hb910b418, 32'hbaa1dfb9, 32'hb8dc3372, 32'h3cd0a88f, 32'hb816feb5, 32'hb816feb5, 32'hbc8e9d52, 32'hb816feb5, 32'h3ede4884, 32'hbed55561, 32'hbf555550, 32'hbed55561, 32'h3fa4a287, 32'hbc441dd2, 32'hbcc41dd2, 32'h3cc41dd2, 32'hbc441dd2, 32'hbc441dd2, 32'h3e088c61, 32'hbd8888b5, 32'hb76ae18b, 32'h3e088ace, 32'hbd8888b5, 32'hb716feb5, 32'h3ced373b, 32'hb58637bd, 32'hb8841ede, 32'hb87fda40, 32'hbcec3116, 32'hbd8888b5, 32'hbd8888b5, 32'h36c9539c, 32'h3eaaacfb, 32'hb80205ff, 32'h36a7c5ac, 32'h358637bd, 32'hbc441dd2, 32'hb76ae18b, 32'hb8a9de8b, 32'h384d8559, 32'h3c684ad8, 32'hbb0ca3e8, 32'hb78e9b39, 32'hbc441dd2, 32'hb716feb5, 32'hb855e8d5, 32'hb88a697b, 32'hbb08722a, 32'h3c689eba, 32'hb7a7c5ac, 32'hb716feb5, 32'hb851b717, 32'hbb09a027, 32'hb88a697b, 32'hb7a7c5ac, 32'hbc441dd2, 32'h3c68ea3a, 32'hbf555550, 32'hbcec3116, 32'hb796feb5, 32'hb796feb5, 32'h3f5cb934, 32'hbf555550, 32'hbed55561, 32'hbc441dd2, 32'hbf555550, 32'h4006df33, 32'hbc441dd2, 32'hb75a1a93, 32'hb80a697b, 32'hb649539c, 32'hb58637bd, 32'hb58637bd, 32'hbcc41dd2, 32'h3cc486ad, 32'hb70637bd, 32'hb7b88ca4, 32'hba61f7d7, 32'hba102de0, 32'h39dbad3a, 32'hbc441dd2, 32'h3c54e4c9, 32'hbd8888b5, 32'h3e088ace, 32'hb716feb5, 32'hbd8888b5, 32'hbd8888b5, 32'hbd8888b5, 32'hbd8888b5, 32'hbe4ccccd, 32'hbc441dd2, 32'hbd8888b5, 32'hbd8888b5, 32'hbe4ccccd, 32'hbcc41dd2, 32'hbd8888b5, 32'h401e86b6, 32'hbd8888b5, 32'hbe4ccccd, 32'hbcc41dd2, 32'hbd8888b5, 32'hbd8888b5, 32'hbe4ccccd, 32'hbcc41dd2, 32'hbd8888b5, 32'hbd8888b5, 32'hbe4ccccd, 32'hbcc41dd2, 32'hbd8888b5, 32'hbd8888b5, 32'hbe4ccccd, 32'hbcc41dd2, 32'hbd8888b5, 32'h3f800000, 32'hbc441dd2, 32'hbe4ccccd, 32'h4170022d, 32'hba017fc7, 32'hb796feb5, 32'hb796feb5, 32'hb58637bd, 32'hba01c2e3, 32'h3b28e2e3, 32'hba8333fd, 32'hba82adc5, 32'hb8ae1049, 32'hb76ae18b, 32'hbc441dd2, 32'hb78637bd, 32'hbaac3a86, 32'h3c518d26, 32'h393fe3b0, 32'h39b2c83f, 32'hbc441dd2, 32'hb716feb5, 32'hb7b88ca4, 32'hba6cb74e, 32'h39ea5b53, 32'h3c558c8f, 32'hba1741d1, 32'hbd8888b5, 32'hbe4ccccd, 32'hbd8888b5, 32'h360637bd, 32'h390d8ec9, 32'hb9755de6, 32'hb969d51b, 32'h3eaad491};
localparam integer A_BRAMInd[0:664] = '{0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 1, 2, 1, 2, 3, 0, 1, 2, 0, 2, 3, 0, 1, 2, 3, 1, 2, 3, 0, 1, 2, 3, 0, 1, 3, 0, 1, 0, 1, 2, 3, 0, 1, 2, 3, 1, 2, 0, 1, 2, 3, 0, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 2, 3, 0, 1, 2, 3, 0, 1, 2, 0, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 0, 1, 3, 3, 0, 1, 2, 0, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 1, 2, 3, 0, 1, 2, 3, 0, 1, 3, 0, 1, 0, 1, 2, 3, 0, 1, 2, 0, 1, 2, 0, 1, 2, 3, 0, 1, 3, 0, 1, 2, 3, 0, 1, 2, 0, 1, 2, 1, 3, 0, 1, 2, 3, 1, 2, 3, 0, 2, 0, 2, 3, 0, 1, 2, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 1, 0, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 1, 2, 1, 2, 0, 3, 0, 1, 0, 1, 3, 0, 1, 2, 2, 3, 0, 1, 2, 3, 1, 3, 1, 0, 2, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 0, 2, 0, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 3, 0, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 0, 1, 2, 3, 0, 1, 3, 0, 1, 2, 3, 0, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 3, 0, 1, 2, 3, 0, 1, 3, 1, 2, 3, 0, 1, 2, 1, 1, 2, 0, 1, 3, 3, 0, 3, 2, 1, 3, 1, 2, 3, 0, 1, 3, 0, 3, 0, 1, 2, 3, 1, 3, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 2, 3, 0, 1, 2, 3, 0, 1, 0, 1, 2, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0, 1, 2, 3, 0};
localparam integer A_BRAMAddr[0:664] = '{0, 0, 0, 0, 1, 1, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 4, 4, 4, 4, 5, 5, 5, 5, 6, 6, 6, 6, 7, 7, 7, 7, 8, 8, 8, 8, 9, 9, 9, 9, 10, 10, 10, 10, 11, 11, 11, 11, 12, 12, 12, 12, 13, 13, 13, 13, 14, 14, 14, 14, 15, 15, 15, 15, 16, 16, 16, 16, 17, 17, 17, 17, 18, 18, 18, 18, 19, 19, 19, 19, 20, 20, 20, 20, 21, 21, 21, 21, 22, 22, 22, 22, 23, 23, 23, 23, 24, 24, 24, 25, 25, 25, 25, 26, 26, 26, 26, 27, 27, 27, 27, 28, 28, 28, 28, 29, 29, 29, 29, 30, 30, 30, 30, 31, 31, 31, 31, 32, 32, 32, 32, 33, 33, 33, 33, 34, 34, 34, 35, 35, 36, 36, 36, 37, 37, 37, 38, 38, 38, 39, 39, 39, 39, 40, 40, 40, 41, 41, 41, 41, 42, 42, 42, 43, 43, 44, 44, 44, 44, 45, 45, 45, 45, 46, 46, 47, 47, 47, 47, 48, 48, 48, 49, 49, 49, 49, 50, 50, 50, 50, 51, 51, 51, 51, 52, 52, 52, 52, 53, 53, 53, 53, 54, 54, 54, 54, 55, 55, 55, 55, 56, 56, 56, 56, 57, 57, 57, 57, 58, 58, 58, 59, 59, 59, 59, 60, 60, 60, 61, 61, 61, 62, 62, 62, 62, 63, 63, 63, 63, 64, 64, 64, 65, 65, 65, 66, 67, 67, 67, 68, 68, 69, 69, 69, 69, 70, 70, 70, 70, 71, 71, 71, 71, 72, 72, 72, 72, 73, 73, 73, 73, 74, 74, 74, 74, 75, 75, 75, 75, 76, 76, 76, 77, 77, 77, 77, 78, 78, 78, 79, 79, 80, 80, 80, 80, 81, 81, 81, 82, 82, 82, 83, 83, 83, 83, 84, 84, 84, 85, 85, 85, 85, 86, 86, 86, 87, 87, 87, 88, 88, 89, 89, 89, 89, 90, 90, 90, 91, 91, 92, 92, 92, 93, 93, 93, 94, 94, 94, 95, 95, 95, 95, 96, 96, 96, 96, 97, 97, 97, 97, 98, 98, 98, 98, 99, 99, 99, 99, 100, 100, 100, 100, 101, 101, 101, 101, 102, 102, 102, 102, 103, 103, 103, 103, 104, 105, 105, 105, 106, 106, 106, 106, 107, 107, 107, 107, 108, 108, 109, 109, 109, 109, 110, 110, 110, 110, 111, 111, 111, 112, 112, 113, 113, 114, 114, 115, 115, 116, 116, 116, 117, 117, 117, 118, 118, 119, 119, 119, 119, 120, 120, 121, 122, 122, 123, 123, 124, 124, 124, 124, 125, 125, 125, 125, 126, 126, 126, 126, 127, 127, 127, 127, 128, 128, 128, 128, 129, 129, 129, 129, 130, 130, 130, 131, 131, 131, 131, 132, 132, 132, 132, 133, 133, 133, 133, 134, 134, 134, 135, 135, 136, 136, 136, 137, 137, 137, 137, 138, 138, 138, 138, 139, 139, 139, 139, 140, 140, 141, 141, 142, 142, 142, 142, 143, 143, 143, 143, 144, 144, 144, 144, 145, 145, 145, 145, 146, 146, 146, 146, 147, 147, 147, 147, 148, 148, 148, 149, 149, 149, 149, 150, 150, 150, 151, 151, 151, 151, 152, 152, 153, 153, 153, 153, 154, 154, 154, 154, 155, 155, 155, 155, 156, 156, 156, 156, 157, 157, 157, 157, 158, 158, 158, 158, 159, 159, 159, 159, 160, 160, 160, 161, 161, 161, 161, 162, 162, 162, 163, 163, 163, 164, 164, 164, 165, 166, 166, 167, 167, 167, 168, 169, 169, 170, 171, 171, 172, 172, 172, 173, 173, 173, 175, 175, 176, 176, 176, 176, 177, 177, 178, 178, 178, 179, 179, 179, 179, 180, 180, 180, 180, 181, 181, 181, 181, 182, 182, 182, 183, 184, 184, 184, 185, 185, 186, 186, 188, 188, 189, 189, 192, 192, 192, 193, 193, 193, 193, 194, 194, 194, 194, 195, 195, 195, 195, 196, 196, 196, 196, 197, 197, 197, 198, 199, 199, 199, 199, 200, 200, 200, 200, 201, 201, 201, 201, 202};

//Constant array to load the instruction BRAM
localparam integer total_instructions = 1268;
localparam integer sub_instructions = 3;
localparam integer Inst[0:1267][0:2] = '{{32'h80000000, 32'h7021010, 32'h6d0},{32'hb0058106, 32'h94421021, 32'h850},{32'h80028000, 32'h4282140e, 32'h670},{32'h90046054, 32'h4703d623, 32'h8e0},{32'hc0034000, 32'h47828418, 32'h8f0},{32'hc0035600, 32'h6d41780b, 32'hff8},{32'h60058000, 32'hb02380c, 32'h8e0},{32'h50044286, 32'h7a423c21, 32'h8f0},{32'ha0044000, 32'h4282d010, 32'h500},{32'hb0056108, 32'h8fc1781e, 32'h5f0},{32'h20028000, 32'hd021803, 32'h860},{32'h9463a502, 32'h76c09010, 32'he48},{32'he0000600, 32'h78c17c0b, 32'h858},{32'h70058012, 32'h7682161c, 32'h850},{32'h86b00080, 32'h4741ac17, 32'hbd0},{32'haa501090, 32'h47c3aa02, 32'h1138},{32'hd0000282, 32'h81421c0b, 32'he40},{32'h28b00010, 32'h47023a12, 32'h920},{32'hcad00010, 32'h4e023e09, 32'h9c0},{32'hb0035402, 32'h30818010, 32'h11d8},{32'h28580400, 32'h49023812, 32'h5f8},{32'h5b180092, 32'hd43ce1e, 32'h850},{32'h60000100, 32'h92c21a10, 32'h840},{32'hf002a002, 32'h92821c0b, 32'h880},{32'h68d00000, 32'h4302181c, 32'h40},{32'hd7600130, 32'h81c38610, 32'h490},{32'h30000004, 32'h4d826c21, 32'hbd8},{32'h80046000, 32'h47024017, 32'h900},{32'hf4e00280, 32'h67444a10, 32'h650},{32'h600000a0, 32'h4e449618, 32'h928},{32'ha0001400, 32'h28838410, 32'h1058},{32'h19700006, 32'h30c27022, 32'h9c0},{32'h40044000, 32'h4942500d, 32'h6b0},{32'h2872a480, 32'h87c06803, 32'h848},{32'h6004a000, 32'h61021411, 32'h8c0},{32'h3b100056, 32'h27043a1e, 32'h888},{32'h20000c00, 32'h50821a14, 32'h11c8},{32'h66680c10, 32'h42026e10, 32'h1048},{32'hc003a000, 32'h23821810, 32'h920},{32'h58d00, 32'h6fc24204, 32'h10d8},{32'h280, 32'h91c21819, 32'h870},{32'ha0028280, 32'h65421801, 32'h570},{32'h30009414, 32'h64027220, 32'h1288},{32'hf0000486, 32'h90407c1f, 32'h6b8},{32'h90000210, 32'h79c06a12, 32'h430},{32'ha0000020, 32'h2b83c20f, 32'h7e0},{32'ha002a030, 32'h78441a01, 32'h8c8},{32'hc0000050, 32'h35040e0e, 32'h6a0},{32'h30035480, 32'h42417014, 32'h1158},{32'hd0001002, 32'hd806c10, 32'h1018},{32'he0046000, 32'h3e01f010, 32'h8c0},{32'h6a746420, 32'h1d843e07, 32'h878},{32'hc0056080, 32'h43c44810, 32'h880},{32'hc9500000, 32'h44809410, 32'h890},{32'h15580028, 32'h7803821f, 32'h870},{32'h6b00000, 32'h3f81fc06, 32'h310},{32'ha662a430, 32'h3f03960f, 32'h7e8},{32'h8003a000, 32'h3e01ac0f, 32'h6c0},{32'hc8556090, 32'h35447210, 32'h8c0},{32'h85700000, 32'hd005003, 32'h1c0},{32'hd4e80018, 32'h2a806e20, 32'h550},{32'h10034012, 32'h3e81f21d, 32'h7d0},{32'h70034402, 32'h44415807, 32'h1118},{32'h80000200, 32'h90c22016, 32'h5d0},{32'h10040284, 32'h8ac12423, 32'h888},{32'hd0001000, 32'h44c1001f, 32'h10b8},{32'ha0000600, 32'h8bc23205, 32'h318},{32'h40001480, 32'h3f41fe0b, 32'h1008},{32'h90000282, 32'h7e42680f, 32'h9b0},{32'h28000, 32'h43844811, 32'h6c8},{32'ha8e80000, 32'h4641f80f, 32'hf08},{32'h9004a090, 32'h2ac3da03, 32'h5b0},{32'h70000084, 32'h3ec0f41f, 32'h3e0},{32'h20028000, 32'h44817c11, 32'h600},{32'h66a8010, 32'h4402220c, 32'h880},{32'h34280, 32'h8d423812, 32'h900},{32'he5280000, 32'h4a83a808, 32'h950},{32'h85180150, 32'h8e444213, 32'h9c0},{32'ha0054000, 32'h4f027013, 32'h100},{32'h6b180420, 32'h29842a0a, 32'h9b8},{32'h40056000, 32'h45022011, 32'h880},{32'hb7284016, 32'h1e01fa22, 32'h1110},{32'he6b00000, 32'h1f813007, 32'h4d0},{32'h266a8400, 32'h8d02b00c, 32'h3e8},{32'hc6680600, 32'h71c2241f, 32'h608},{32'h3a600080, 32'h4441bc11, 32'h6b0},{32'ha8b01000, 32'h44022822, 32'h12a8},{32'h1ae00000, 32'h50027c12, 32'h140},{32'h98580022, 32'h4ac43613, 32'h60},{32'h90000004, 32'h1d80ec1f, 32'h540},{32'h74746002, 32'h4f44700a, 32'h720},{32'h15300002, 32'h44023011, 32'hf00},{32'h54e00000, 32'h8f814011, 32'he0},{32'h96600500, 32'h86c01c07, 32'h4d8},{32'hf0001000, 32'h29814c07, 32'hfa8},{32'h30046000, 32'h4383800c, 32'h8a0},{32'h8d00000, 32'h45022611, 32'h8b0},{32'hf7500000, 32'h9541a80d, 32'h6a0},{32'h60044000, 32'h90022a0d, 32'h6c0},{32'hcad00000, 32'h5041800b, 32'h610},{32'h99500012, 32'h980ee22, 32'h130},{32'ha0034000, 32'h4e015213, 32'h9e0},{32'head01450, 32'h39442601, 32'hdc8},{32'h1400, 32'h18823206, 32'h10a8},{32'h3a000, 32'h2a01420f, 32'h540},{32'h24580290, 32'h74c14e06, 32'h320},{32'h2a000, 32'h44804c11, 32'h130},{32'h47444000, 32'h49826813, 32'h1130},{32'hd4758016, 32'h4101aa1b, 32'h8b8},{32'h40000c00, 32'h3600b405, 32'hea8},{32'h10030058, 32'h62048624, 32'h6c8},{32'hd0000086, 32'h9c03022, 32'h618},{32'h80001000, 32'h46022011, 32'hf58},{32'h47280000, 32'h600cc06, 32'h9e8},{32'haa600c80, 32'h18c0f407, 32'hf98},{32'h40058000, 32'h19815006, 32'h310},{32'h4a9c0400, 32'h2a40e807, 32'h328},{32'he0058010, 32'h8d004e0b, 32'h610},{32'h57500012, 32'h2c036a13, 32'h8a8},{32'h90000030, 32'h1f048a0d, 32'h3f0},{32'h70026082, 32'h3641f423, 32'h7d0},{32'h60044000, 32'h87822c16, 32'h8d0},{32'h8d00280, 32'h66c1fc1d, 32'h7f0},{32'h45600000, 32'h4e807013, 32'h9e0},{32'h97500230, 32'h82c36e11, 32'h410},{32'hb4700102, 32'h8940ce07, 32'h1c0},{32'hf0000414, 32'h17815220, 32'h1228},{32'h50000032, 32'h19c3ca07, 32'h9f0},{32'hc0000020, 32'h30836209, 32'h4d0},{32'h8ab30000, 32'h82806c03, 32'h618},{32'h77280418, 32'h1b83c61e, 32'h3f8},{32'h30000016, 32'h2301f622, 32'h470},{32'ha0026000, 32'h23043810, 32'h10d0},{32'hc9426000, 32'h3101880b, 32'h330},{32'h77600004, 32'h3f01fe1d, 32'hea0},{32'ha4f00000, 32'h1f80fc07, 32'h9e8},{32'h67600000, 32'h36810623, 32'h6d0},{32'h45580000, 32'h1c80f007, 32'h3c0},{32'h756002a6, 32'h8c446222, 32'h740},{32'h200000a0, 32'h30c3d213, 32'h9a0},{32'hc002a000, 32'he813e0f, 32'h2b0},{32'h90030150, 32'h77439a03, 32'h2c0},{32'hb0000484, 32'h7ac1441d, 32'h478},{32'h70001082, 32'h23c29825, 32'h1298},{32'ha0000200, 32'h6bc3980f, 32'h8d8},{32'h4004a000, 32'h31018a0c, 32'h5f0},{32'h56a80000, 32'h8b80ec10, 32'h400},{32'h67320000, 32'h1980fe1d, 32'h320},{32'hea980000, 32'h36c06820, 32'h1d0},{32'h2b100200, 32'h77c0f20c, 32'h610},{32'h50054402, 32'h1f00f81b, 32'h9a8},{32'h46080, 32'hec18415, 32'h610},{32'h60044050, 32'h4d835a13, 32'hc90},{32'h40056120, 32'h65c46e09, 32'h4b0},{32'ha002a000, 32'h4003940a, 32'h560},{32'hd85aa002, 32'h43843c0f, 32'h8d0},{32'h88d00000, 32'h3081880d, 32'h6c0},{32'hf8c54432, 32'h203461c, 32'h408},{32'h10000030, 32'h88c40208, 32'hc70},{32'h80000020, 32'h19c3fa03, 32'h4f0},{32'h3000a112, 32'h8f43ae0c, 32'h810},{32'h20000510, 32'h72c0fa15, 32'h1188},{32'h80000290, 32'h8b418608, 32'h450},{32'h7002a002, 32'h2700e813, 32'h3b0},{32'h66728400, 32'h90815c0a, 32'h4b8},{32'he7600400, 32'h3601fc0d, 32'h568},{32'haf08000, 32'h46015411, 32'h550},{32'h97444012, 32'h2c04aa0d, 32'h560},{32'h56b00000, 32'h4f036c0c, 32'h9b0},{32'he8980020, 32'h3283660b, 32'h650},{32'h85580400, 32'h1e00f022, 32'h1d8},{32'ha7600000, 32'hf03cc03, 32'h810},{32'hcb180020, 32'h1f03e607, 32'h890},{32'hb0056484, 32'h7bc4601f, 32'h458},{32'he8700400, 32'h4f836813, 32'h3b8},{32'he7280000, 32'h2a813a15, 32'h570},{32'h54c01492, 32'h40447a1d, 32'h10f8},{32'h20000010, 32'h95c15617, 32'h708},{32'he0000280, 32'h73c0fc07, 32'h8d8},{32'h40058000, 32'h3581620d, 32'h980},{32'h9003a004, 32'h4f42901b, 32'h9a0},{32'hb8b00000, 32'h32c30824, 32'h3d0},{32'h40021000, 32'h2580f209, 32'hcd8},{32'hd003a402, 32'hf405c07, 32'h1128},{32'h10000008, 32'h2180f020, 32'h1120},{32'hc6b08000, 32'h4e027c04, 32'h270},{32'ha8c2a200, 32'h6dc2241f, 32'h870},{32'haaa00000, 32'h2b015e0a, 32'hc00},{32'h4003a100, 32'h6643601b, 32'ha00},{32'hf9500402, 32'h23011807, 32'he88},{32'h80046080, 32'h35c0f007, 32'h9d0},{32'h80058100, 32'h6e427813, 32'hdc0},{32'h95600480, 32'h7dc12c14, 32'h3d8},{32'hb8700082, 32'h25c1e823, 32'he80},{32'h8b01000, 32'h4082001d, 32'h11b8},{32'h39580482, 32'h1ec18423, 32'h1198},{32'h70000600, 32'h68c20008, 32'h278},{32'hf0000200, 32'h83c35e13, 32'h8a0},{32'h60020080, 32'h2b422602, 32'h130},{32'h60054000, 32'h4f836400, 32'h30},{32'h67054010, 32'h30811a0c, 32'h640},{32'h9ad00012, 32'h15044607, 32'h270},{32'h66b00030, 32'h3584820d, 32'ha10},{32'haf00100, 32'h6cc27a08, 32'h1190},{32'heab00000, 32'h5981e81c, 32'h4c8},{32'h59700c00, 32'h3681b40f, 32'h1168},{32'h20046000, 32'h40c22411, 32'hb80},{32'h30058004, 32'h4202501a, 32'h960},{32'h88d00480, 32'h71413009, 32'h8a8},{32'h70058002, 32'h2027402, 32'h50},{32'h76501082, 32'h69c01400, 32'hdb8},{32'h50000008, 32'h90814c1f, 32'ha08},{32'h87300000, 32'h22848e08, 32'h648},{32'h3a000, 32'h7d80aa08, 32'h6c0},{32'h8af04000, 32'h71022814, 32'h8b0},{32'h28d01400, 32'h21404402, 32'hd98},{32'h30058012, 32'h5181b624, 32'h7b8},{32'h30000c32, 32'h2043211, 32'h11e8},{32'h70000006, 32'h8e023c24, 32'h600},{32'h97000102, 32'h93406409, 32'h190},{32'h80044000, 32'h7102300f, 32'h8d0},{32'h48d00280, 32'h75c18c0c, 32'h58},{32'h2004a000, 32'h1980cc21, 32'h4a0},{32'hda546480, 32'h22c4060a, 32'h1108},{32'h20000090, 32'h94c1b223, 32'h430},{32'h5700000, 32'h81005800, 32'h428},{32'h36600002, 32'h2b041802, 32'h8b8},{32'h28f00000, 32'h4083e411, 32'h7e0},{32'ha8981400, 32'h77807803, 32'he38},{32'hcae00000, 32'h2302f008, 32'h220},{32'h14756018, 32'h3c80661a, 32'h968},{32'h30000006, 32'h6d82701d, 32'ha00},{32'h27100010, 32'h4d018e13, 32'h8d8},{32'h6003a410, 32'hd80ce03, 32'he58},{32'h20056000, 32'h4e028414, 32'h4a8},{32'h48e80000, 32'h48022811, 32'he30},{32'h18a80006, 32'h2240441c, 32'h120},{32'he0028000, 32'h75805a0f, 32'h7f0},{32'hf4e80000, 32'h2081040a, 32'h1180},{32'h96a00000, 32'h40c2d41c, 32'h740},{32'hd4701002, 32'h4a807a08, 32'hef8},{32'h70000030, 32'h6e047604, 32'h9c0},{32'h34000, 32'h26813400, 32'h9f0},{32'hf4746082, 32'h4d42a823, 32'ha08},{32'h70001002, 32'h4e029803, 32'hd88},{32'h28f00000, 32'h6d027002, 32'ha20},{32'h37101400, 32'h84400014, 32'hed8},{32'h50000400, 32'h8c01d411, 32'h128},{32'h48f00000, 32'h3f039411, 32'h8b0},{32'h28c2a000, 32'h42010008, 32'h1110},{32'h48a80c00, 32'h45810611, 32'he28},{32'h6003a000, 32'h1981d206, 32'h3d0},{32'h10056404, 32'h2000fc1e, 32'h9d8},{32'ha0038010, 32'h27813623, 32'h11c0},{32'h85580000, 32'ha028202, 32'hed0},{32'h6a80000, 32'h6b827000, 32'ha70},{32'hd7100000, 32'h82422c14, 32'he20},{32'h8b00000, 32'h4782401c, 32'ha28},{32'h8ae00000, 32'h2680001b, 32'h4e0},{32'hba726400, 32'h7b41fc0e, 32'h8b8},{32'h40008000, 32'h88844400, 32'h20},{32'ha7054080, 32'h45c0d80e, 32'h360},{32'h74601402, 32'h9504a806, 32'h12b8},{32'h87300080, 32'h20423011, 32'he30},{32'h88a80000, 32'h1480a409, 32'h11d0},{32'h25446000, 32'h9805000, 32'h10},{32'h8c54000, 32'h48823c1c, 32'h8b0},{32'hab180100, 32'h88411408, 32'ha78},{32'h58000, 32'h46c13412, 32'h1290},{32'h25350400, 32'h19024206, 32'h4e8},{32'hf003a002, 32'h4c42400f, 32'h910},{32'h50028012, 32'h89033600, 32'h3e0},{32'he6800000, 32'hf00780f, 32'h1d0},{32'h96a00e86, 32'h8340da1e, 32'h1078},{32'h10000000, 32'h4584340e, 32'h130},{32'h90f44010, 32'h8f00a611, 32'h4e0},{32'h36b00402, 32'h27c2cc00, 32'hec8},{32'h90001000, 32'h39024002, 32'hd28},{32'hb0008c02, 32'h49824c08, 32'h1258},{32'h16600002, 32'h68818812, 32'h630},{32'h38d00480, 32'h1942740a, 32'h1148},{32'h70000408, 32'h900481b, 32'h918},{32'h46000, 32'h2080a005, 32'h1120},{32'h6858000, 32'h4a825412, 32'h1f0},{32'h47620000, 32'hb807a21, 32'h120},{32'hba580484, 32'h7c428c20, 32'h148},{32'h30000008, 32'h3602361b, 32'h1250},{32'hf4f00000, 32'h67023c09, 32'h0},{32'h67300080, 32'h48c26c1b, 32'h9e0},{32'h6b100000, 32'h49810412, 32'h910},{32'h46a81000, 32'h4c024e0c, 32'hf18},{32'hb000a006, 32'h1200001b, 32'h250},{32'h66500010, 32'h16004a06, 32'h2c0},{32'h14581402, 32'h5802c05, 32'hd18},{32'h30046400, 32'h4802408, 32'h1f8},{32'h46000, 32'h49025612, 32'h920},{32'h65580000, 32'hbc27813, 32'hdb0},{32'h5600000, 32'h3901b000, 32'h730},{32'ha7100000, 32'h2681ca09, 32'hf88},{32'hb0056000, 32'h4f000017, 32'h1f0},{32'hd0030004, 32'h500281e, 32'h9e8},{32'h70046400, 32'h60830412, 32'h638},{32'h46000, 32'h78804c00, 32'h0},{32'h87054000, 32'h2e817401, 32'hf50},{32'h46c6410, 32'h16402e00, 32'h11a8},{32'hc0000410, 32'h13802604, 32'h1098},{32'h2003a000, 32'h3181880c, 32'h930},{32'h495a0000, 32'h4941500b, 32'h9e0},{32'h8b304000, 32'h2a01440a, 32'h520},{32'hb8556002, 32'h66833409, 32'h738},{32'hc7300080, 32'h4f402401, 32'h1280},{32'h45280010, 32'h2a18, 32'hcd0},{32'h94680012, 32'h62830619, 32'h1050},{32'h14580002, 32'h6f824800, 32'h910},{32'h86a00010, 32'h7b017607, 32'h258},{32'h97700000, 32'hc809c01, 32'h190},{32'hc8734480, 32'h13c25c12, 32'h1218},{32'h4a600410, 32'h4220c, 32'h938},{32'ha010, 32'h7e027a00, 32'h5c0},{32'h96500002, 32'h2dc00c0a, 32'h30},{32'he0044000, 32'h50027813, 32'h528},{32'hfb180000, 32'h2817, 32'he0},{32'h45000000, 32'h48800012, 32'h920},{32'h54e80000, 32'h48847418, 32'h960},{32'h88d00000, 32'h62c0d006, 32'h310},{32'h88a80000, 32'h88024a11, 32'h8d0},{32'h3ad00080, 32'hcc00025, 32'h768},{32'h20000000, 32'h7a01900c, 32'h288},{32'ha7600080, 32'h31c25e0e, 32'h3d0},{32'h6ab00000, 32'h1481541f, 32'h2a0},{32'h7b026012, 32'h20000e1a, 32'hf10},{32'hc4f00000, 32'h4880001b, 32'h940},{32'h6ad00000, 32'h50412c09, 32'h4b0},{32'hd8a80000, 32'h49024801, 32'h0},{32'h50046000, 32'h4a024c12, 32'h930},{32'h48980000, 32'h49000012, 32'h968},{32'h90056000, 32'h46800006, 32'h0},{32'h80030000, 32'h8382040f, 32'h8d8},{32'h47600000, 32'h3182c816, 32'h640},{32'h4c58000, 32'h77011400, 32'h460},{32'h86728400, 32'h3b44040a, 32'h2a8},{32'ha9700000, 32'h30819424, 32'h5c8},{32'haae00000, 32'h4a810a12, 32'h910},{32'h6a80000, 32'h26004c20, 32'h948},{32'h7b330410, 32'h24a09, 32'hd08},{32'h60000000, 32'h24c12, 32'hd00},{32'h58a80012, 32'h4a433e12, 32'h0},{32'h40000080, 32'h46c24c12, 32'h940},{32'h9500000, 32'h3e823410, 32'h8d0},{32'h5ac44012, 32'h1832a16, 32'h30},{32'ha0034400, 32'h4681921b, 32'h468},{32'h7af00000, 32'h4b025405, 32'h930},{32'ha8980000, 32'h3281840c, 32'h588},{32'h27280000, 32'h1901961a, 32'hfb8},{32'hbaf00090, 32'h26444e12, 32'h0},{32'hc0000000, 32'h4b833c12, 32'h188},{32'hab180000, 32'h25412, 32'hd00},{32'h78a80000, 32'h7b811c12, 32'h480},{32'h88d00000, 32'h4580001b, 32'h990},{32'had00090, 32'h6f423600, 32'h948},{32'h60000080, 32'h1c20612, 32'h940},{32'h8002a000, 32'h46800012, 32'h960},{32'h6ad00000, 32'h6ec26203, 32'hb60},{32'h5700000, 32'h4b419400, 32'h630},{32'h68800000, 32'h4a032812, 32'hc00},{32'h8533a000, 32'h6f000012, 32'hb98},{32'hcaf00000, 32'h1824812, 32'h970},{32'hb100030, 32'h4bc37a00, 32'h0},{32'hb0000000, 32'h3f81f812, 32'h800},{32'h7100000, 32'h4c023400, 32'h488},{32'he7000000, 32'h4f000013, 32'ha00},{32'haad00480, 32'h8ec0a405, 32'h948},{32'h4b300000, 32'h5825412, 32'hf90},{32'hc9426000, 32'h15c0a, 32'h1220},{32'heaa00000, 32'h5bc11808, 32'h480},{32'hbb100480, 32'h4a43ee0c, 32'hdf8},{32'h10000000, 32'h41020818, 32'h7e0},{32'ha6a00000, 32'h4b025a12, 32'hdf0},{32'h2a980000, 32'h1483b605, 32'h978},{32'h20056000, 32'h4f01fc14, 32'ha20},{32'had08000, 32'h4b83b400, 32'h940},{32'h8980000, 32'h28000, 32'h998},{32'ha0040000, 32'h3c21, 32'ha08},{32'ha600090, 32'h6442e00, 32'h2e8},{32'h20000000, 32'h3701b824, 32'h968},{32'ha7600000, 32'h8e815e12, 32'h960},{32'h6ad00000, 32'h3201840c, 32'h488},{32'hb180000, 32'h4101f800, 32'h830},{32'h67100000, 32'h5820a01, 32'h2b0},{32'h34756002, 32'h4b40a005, 32'h290},{32'he0028480, 32'h7240bc05, 32'h808},{32'h60058000, 32'h82807403, 32'ha28},{32'h7600010, 32'h4bc28200, 32'hde8},{32'h0, 32'h2b815c00, 32'h560},{32'h6a00000, 32'h50003e00, 32'ha00},{32'h20034000, 32'h37810408, 32'he80},{32'h8ab0000, 32'h4b01ba00, 32'h0},{32'h30000, 32'h2b04880b, 32'h968},{32'h8e80000, 32'h32403000, 32'hd0},{32'h78500012, 32'h49e01, 32'h838},{32'h40000400, 32'h900ae02, 32'h298},{32'hf0056002, 32'h25805, 32'h960},{32'h80044000, 32'h3f020403, 32'h810},{32'hc4e0a000, 32'he828003, 32'h1070},{32'h84e80200, 32'h6b400414, 32'h10},{32'h2a744080, 32'h50415e1d, 32'h7a0},{32'ha500080, 32'h37c26013, 32'h0},{32'h38680080, 32'h4b400008, 32'h0},{32'he0044000, 32'h50007c03, 32'h1d0},{32'h18a80030, 32'h6b04160b, 32'ha20},{32'he4f00000, 32'h15c0a, 32'hd8},{32'h50058002, 32'h21810c02, 32'h1180},{32'h86a00010, 32'hf825a1e, 32'h0},{32'hea580410, 32'h4080760f, 32'hf48},{32'h7400000, 32'h5a007800, 32'hd20},{32'h64588090, 32'h7d400609, 32'h4c0},{32'h2002a000, 32'h6c410808, 32'ha58},{32'he004a000, 32'h4b825812, 32'h7a8},{32'h17280010, 32'h5800213, 32'hc0},{32'h26000, 32'h10000013, 32'h1f0},{32'hf0980050, 32'h80437603, 32'h0},{32'hf0000082, 32'h91428a0a, 32'h0},{32'h0, 32'h3c01e, 32'h440},{32'h29500000, 32'h21010e08, 32'hf68},{32'ha003a000, 32'hfc1b00d, 32'h6d0},{32'hd5280402, 32'h20603, 32'hdd8},{32'h20000400, 32'h5a400025, 32'h4c8},{32'h5a700418, 32'h10a19, 32'hf78},{32'h80000000, 32'h6803001, 32'hd0},{32'hf85aa400, 32'hc809412, 32'hc8},{32'h68f00000, 32'h28c14, 32'h7e0},{32'h28a80000, 32'h1041f810, 32'h810},{32'h5280000, 32'h1880d000, 32'h350},{32'h8d00000, 32'h2183c400, 32'hc0},{32'h77000484, 32'h21400020, 32'he78},{32'h60000000, 32'h36844408, 32'h430},{32'h5286000, 32'h32048c00, 32'h630},{32'h8980000, 32'h27813800, 32'h4c0},{32'h8980000, 32'h9101600b, 32'h788},{32'h88e80410, 32'h3de01, 32'hd8},{32'ha000, 32'h4a025c00, 32'h970},{32'hb4e00000, 32'h2003e204, 32'hf60},{32'h74f00000, 32'h40800014, 32'h800},{32'h86800000, 32'h500cc06, 32'hb0},{32'heb026000, 32'h810c1c, 32'h10},{32'h9434000, 32'h3581c000, 32'h12a0},{32'hb4e00012, 32'h104a60d, 32'h20},{32'h70034000, 32'h73819008, 32'h600},{32'h6b40000, 32'h32413400, 32'h4f0},{32'h65000000, 32'h1100881e, 32'h590},{32'h17620480, 32'h6c0000b, 32'hd68},{32'h0, 32'h4b000000, 32'hde0},{32'h4c00000, 32'h6e825800, 32'h990},{32'h87100000, 32'h11216, 32'h0},{32'h3a734410, 32'h34e10, 32'hb8},{32'hd0000082, 32'hc00021, 32'h358},{32'he0000000, 32'h9480000d, 32'h448},{32'h2ac00080, 32'h1420410, 32'h0},{32'hf0058012, 32'h8181921e, 32'h30},{32'h50034000, 32'h24011c17, 32'h1100},{32'h8980400, 32'h27c00000, 32'h598},{32'hd0000000, 32'h60808a24, 32'hc20},{32'he0026000, 32'h2083c412, 32'h420},{32'ha7150000, 32'h25e16, 32'h1160},{32'h4680080, 32'h400000, 32'h998},{32'h20000000, 32'h7b82fe09, 32'h490},{32'h44e80000, 32'h83020810, 32'h0},{32'ha8e80000, 32'hf80780d, 32'h700},{32'h35438002, 32'h2840010, 32'h0},{32'h8580480, 32'h7cc00000, 32'h48},{32'hc0000000, 32'h4844008, 32'ha0},{32'ha9426000, 32'h61830806, 32'h350},{32'h785d4402, 32'he808819, 32'hc28},{32'hf8f00002, 32'h3801b412, 32'h700},{32'hc5180000, 32'h3704a40d, 32'h428},{32'hb7280000, 32'he807c16, 32'h200},{32'h28d00000, 32'h4811801, 32'h10b0},{32'hc5056000, 32'h4180000f, 32'hea0},{32'h55580480, 32'hfc39210, 32'he08},{32'h60000000, 32'h5101c213, 32'h1040},{32'he5580000, 32'h2c37412, 32'h990},{32'h9500480, 32'h86400000, 32'ha8},{32'hb0000002, 32'h24408806, 32'h1d0},{32'h68b00000, 32'h61c10c08, 32'he80},{32'h48a80000, 32'h9805821, 32'h238},{32'h5ae00000, 32'h3841b825, 32'h0},{32'hc0008000, 32'h80000803, 32'h20},{32'h37444082, 32'h85400001, 32'h0},{32'h30000000, 32'h9, 32'h10c8},{32'he0000000, 32'h41c1041c, 32'h420},{32'h89500000, 32'h24028413, 32'h480},{32'h69434000, 32'h1902641d, 32'h340},{32'had40000, 32'h23844009, 32'h998},{32'h8e80000, 32'h11800000, 32'h1f0},{32'h50980000, 32'h85c2c804, 32'hb30},{32'h70028000, 32'h3c80bc08, 32'h300},{32'hd6728002, 32'h4c805a0d, 32'h990},{32'h40034010, 32'h10000a0f, 32'he70},{32'hcab30000, 32'h3801c00d, 32'h208},{32'hc7600000, 32'h42413, 32'h9d0},{32'h28a80000, 32'h1b80dc08, 32'h320},{32'h26a0a090, 32'h24445603, 32'h1a0},{32'h3002a012, 32'h5142661c, 32'h0},{32'h20000000, 32'h51027814, 32'h348},{32'h1b180000, 32'h19805809, 32'h340},{32'h50026418, 32'h11c33223, 32'hb38},{32'ha0000400, 32'h15, 32'h308},{32'h9a700082, 32'h4cc1e620, 32'h0},{32'h90, 32'h10440a09, 32'h480},{32'ha0054000, 32'h3dc13c09, 32'h4f0},{32'h45600000, 32'h3781c225, 32'h9e0},{32'heaf04480, 32'h74400815, 32'h428},{32'h2b300400, 32'h6080de18, 32'h1a8},{32'h80056000, 32'h9400000d, 32'h6e0},{32'h87500000, 32'h3881c020, 32'ha10},{32'h45438410, 32'h5038a01, 32'h348},{32'h80056000, 32'h28000009, 32'h500},{32'h5580000, 32'h3e843000, 32'ha40},{32'h8d00000, 32'h6ac00000, 32'hae8},{32'h10000012, 32'h4ae09, 32'h1a0},{32'h20, 32'h2784a200, 32'h0},{32'hd0006402, 32'h1c013, 32'hda8},{32'h20008000, 32'h6083081e, 32'hc30},{32'h38556002, 32'h6c826418, 32'hb18},{32'h7300000, 32'h1f410, 32'h820},{32'h2b100080, 32'h38c00018, 32'h6e8},{32'h50001402, 32'h51400001, 32'h1068},{32'h40000000, 32'h51041401, 32'ha20},{32'h5181400, 32'h28400000, 32'h1178},{32'h20000000, 32'h5201f81b, 32'ha48},{32'hb180000, 32'h36800000, 32'h6e0},{32'h20026410, 32'h13e15, 32'h1208},{32'ha700480, 32'h75400000, 32'h718},{32'h40000090, 32'h61445e18, 32'h0},{32'ha000, 32'h3f028c00, 32'ha40},{32'hc8d00000, 32'h7280000f, 32'ha38},{32'h87400000, 32'h1a800006, 32'hd10},{32'ha980000, 32'h1b00cc00, 32'h360},{32'ha5180000, 32'ha028820, 32'h150},{32'h7540000, 32'h51427c14, 32'h9d0},{32'h68a80000, 32'h14, 32'h800},{32'h1a800402, 32'h38800025, 32'h6e8},{32'h40000c00, 32'h4182081d, 32'hd78},{32'h89580000, 32'h55400018, 32'h1050},{32'he5280400, 32'h26013809, 32'hc38},{32'h68e80000, 32'h83000014, 32'h0},{32'h8ac00000, 32'h4000001c, 32'h0},{32'h6ac00000, 32'ha805002, 32'h350},{32'h9584000, 32'h5281f400, 32'h11e0},{32'h15180012, 32'h1b428a1b, 32'h0},{32'he0000000, 32'h9805c02, 32'h158},{32'h18e80000, 32'h93049414, 32'h660},{32'hc8d00000, 32'h52404c20, 32'h150},{32'hb100000, 32'h1b035c14, 32'hda0},{32'hf8a80006, 32'h41c28821, 32'hae0},{32'h95300000, 32'h2781e418, 32'hd70},{32'h8b06000, 32'h72020800, 32'h830},{32'hd8d00000, 32'h23, 32'ha48},{32'h80000080, 32'h1ac00002, 32'h828},{32'hc000a000, 32'h51028c0f, 32'ha30},{32'h49426000, 32'h56020401, 32'h820},{32'h67728000, 32'hc005c02, 32'h0},{32'hf9580000, 32'h28014002, 32'h1200},{32'h86a00000, 32'h2, 32'h668},{32'he000a000, 32'h1a80d821, 32'ha00},{32'hae04000, 32'h56034c00, 32'haf0},{32'hf7100402, 32'h57400009, 32'h1088},{32'h20000000, 32'h3d439010, 32'h0},{32'h69400000, 32'hb000002, 32'h170},{32'h7500090, 32'hac3be00, 32'h0},{32'h40000410, 32'h61835618, 32'ha38},{32'h3a400, 32'h52c00000, 32'h828},{32'h20000000, 32'h3282b60c, 32'h660},{32'he7500000, 32'hc409c04, 32'h270},{32'h8a80480, 32'h79414200, 32'h158},{32'h10000012, 32'h41214, 32'h0},{32'hc0000000, 32'h4f00da14, 32'ha70},{32'h6ad00000, 32'h52847814, 32'haf8},{32'hab180000, 32'h24820c08, 32'h4a0},{32'h7540000, 32'ha805800, 32'h838},{32'h68c00000, 32'h62000019, 32'hc50},{32'h27500080, 32'h61c15420, 32'h580},{32'hb100000, 32'h3a011800, 32'h740},{32'h5180000, 32'h31819400, 32'h0},{32'h28c00000, 32'h1401640b, 32'h590},{32'hf8ab0000, 32'h2d83d804, 32'h5b0},{32'he5180000, 32'h12008, 32'h470},{32'h8aa00000, 32'h53829813, 32'h0},{32'ha9580000, 32'h3b81d808, 32'ha78},{32'he9580010, 32'h52c20e04, 32'h280},{32'h8002a000, 32'h9809004, 32'h4a8},{32'h8e80000, 32'hf808404, 32'h178},{32'hae00000, 32'h15c00, 32'hc58},{32'h8000, 32'h7a83d000, 32'h750},{32'ha8d00000, 32'h3a41900c, 32'heb8},{32'hcb000080, 32'h14412408, 32'h4a0},{32'h39500000, 32'h7980800b, 32'hf40},{32'hc6a00000, 32'h2dc1180e, 32'h770},{32'hcb100000, 32'h91812203, 32'h210},{32'hc7500000, 32'h53c00008, 32'h1150},{32'h55400402, 32'h6c035424, 32'h288},{32'h67300000, 32'h12809002, 32'h0},{32'h99580000, 32'h2c816004, 32'h0},{32'h8580400, 32'h8600, 32'h588},{32'h0, 32'h12000, 32'h480},{32'h44000, 32'h19800, 32'h758},{32'h20040000, 32'h24000009, 32'h668},{32'heac00000, 32'hf800003, 32'h580},{32'h6ac00020, 32'h7403f208, 32'h440},{32'head00000, 32'h2d816c0a, 32'h778},{32'hc7600000, 32'h53827814, 32'h218},{32'h8b180000, 32'h3bc0d406, 32'h340},{32'h8aa00000, 32'h3bc04, 32'ha68},{32'hb000000, 32'h37000025, 32'h6f0},{32'he7500000, 32'h2cc0dc06, 32'he50},{32'h98a80012, 32'h6b012225, 32'ha70},{32'h4f00090, 32'h93c19a14, 32'hd90},{32'h45700000, 32'h1b40e, 32'hf80},{32'h5280000, 32'h2c80000b, 32'h4a8},{32'h8003a000, 32'h33808223, 32'h630},{32'ha980000, 32'h29044c22, 32'h448},{32'h2b180000, 32'h52016e10, 32'ha40},{32'h5580000, 32'h53c00000, 32'h350},{32'h80004000, 32'h18c0c, 32'h640},{32'h5280000, 32'h12c1b800, 32'h0},{32'h60008000, 32'hdc06, 32'h380},{32'hf9500000, 32'h89c08006, 32'h200},{32'h40044000, 32'h41829e10, 32'h820},{32'ha980000, 32'h37829600, 32'h0},{32'h50f00080, 32'h2cc1400e, 32'h510},{32'h28000, 32'h31819c00, 32'h670},{32'h44e00000, 32'h33c1440e, 32'h4e0},{32'hc8800280, 32'h96438806, 32'h360},{32'h5280010, 32'h5240d600, 32'h11f8},{32'h40000000, 32'h32028414, 32'h9d0},{32'h8a86400, 32'h2c816400, 32'h6f8},{32'he8f00000, 32'h1a800006, 32'h0},{32'hac00090, 32'h7fc08200, 32'h0},{32'he0000000, 32'hc03bc02, 32'h830},{32'hb184000, 32'h3401a400, 32'h0},{32'h26600400, 32'h2d01ce0b, 32'h518},{32'he003a000, 32'h3380001e, 32'h0},{32'h27400000, 32'h2880000a, 32'h4c0},{32'h6a80000, 32'h29416c00, 32'h590},{32'hd8b00000, 32'h33018c06, 32'hfb0},{32'h95180012, 32'h8404660c, 32'hda0},{32'h26800000, 32'h1584800b, 32'h1210},{32'h2898a000, 32'h1c000022, 32'h1140},{32'h5a980000, 32'h2a822, 32'h388},{32'h8700090, 32'h41c47e00, 32'h0},{32'ha0000000, 32'hc41c80d, 32'h730},{32'h9500480, 32'h2d41a600, 32'h1248},{32'he0000000, 32'h18c0c, 32'h670},{32'h5280000, 32'h92419e00, 32'h0},{32'h30000000, 32'h5384140a, 32'ha70},{32'h75180000, 32'h2401d00b, 32'heb0},{32'h4e00000, 32'h33441000, 32'ha20},{32'h5000480, 32'h7ec00000, 32'h5a8},{32'h0, 32'h15c0dc00, 32'h340},{32'h28800000, 32'h55800015, 32'hd70},{32'h5a980000, 32'h1580a815, 32'h280},{32'hc8980000, 32'h9600000d, 32'h0},{32'hc7400000, 32'h85800003, 32'h230},{32'h7500000, 32'h33846400, 32'h0},{32'hc7000000, 32'h52800023, 32'h820},{32'hea980000, 32'h2d029814, 32'h9d0},{32'h8a80030, 32'h53c41e00, 32'h0},{32'h0, 32'h5101d200, 32'h12c8},{32'h6000, 32'h10800004, 32'h1f0},{32'hea980000, 32'h5380d406, 32'h0},{32'hcb000030, 32'h81037e02, 32'h120},{32'h6a80000, 32'h55c48405, 32'h0},{32'h9400000, 32'h3981c400, 32'h1240},{32'h88980000, 32'h3303ec0c, 32'h738},{32'hc9580000, 32'h1b00d406, 32'h238},{32'hf7280000, 32'h47c0c, 32'h11f0},{32'h5000000, 32'h82000000, 32'hda0},{32'h6800000, 32'h0, 32'hae0},{32'h54700402, 32'h92019814, 32'h1028},{32'h7300000, 32'h40800, 32'h210},{32'h25000000, 32'h13c0a, 32'h520},{32'hb100000, 32'h1c404800, 32'h160},{32'h5000000, 32'ha400, 32'h2b0},{32'h5000000, 32'h1a800, 32'h720},{32'h5000000, 32'h2800000a, 32'h1080},{32'h66a80000, 32'h33411008, 32'hf70},{32'hdaa00000, 32'h33000006, 32'h660},{32'h34000, 32'h52c41000, 32'ha70},{32'he5000000, 32'h52829023, 32'h0},{32'h9580000, 32'h9582ba0e, 32'h6e0},{32'h6a80000, 32'h53829c1b, 32'h688},{32'hc7600000, 32'h10c0d806, 32'h0},{32'h60058000, 32'h84c41c0b, 32'h528},{32'hdb300000, 32'h25012402, 32'h470},{32'h88980000, 32'h15c0000d, 32'h1250},{32'h25400000, 32'h3b014025, 32'h420},{32'hca988000, 32'hb004c02, 32'h440},{32'h7284090, 32'h33449a00, 32'h0},{32'h0, 32'h53800000, 32'h1020},{32'h86800000, 32'h28014, 32'h0},{32'hb000000, 32'h38000000, 32'h6f0},{32'h6800000, 32'h37c00, 32'ha30},{32'hd8b00002, 32'h29e06, 32'h1038},{32'hc0000000, 32'h24812806, 32'h460},{32'h26a01400, 32'h2e412009, 32'h12d8},{32'hb000000, 32'h34000000, 32'h0},{32'h16700002, 32'h39c4980a, 32'h690},{32'h5300010, 32'h3b411200, 32'h0},{32'hd0000000, 32'h3b845402, 32'h770},{32'hc5180000, 32'h5802, 32'h150},{32'hf8a80000, 32'h28814, 32'ha50},{32'h65000000, 32'h2201c008, 32'he70},{32'h4a988000, 32'h7400000f, 32'h7b0},{32'h4ad00000, 32'h5440ac05, 32'h290},{32'haa00000, 32'h23811000, 32'h10b0},{32'h4c00200, 32'h8dc00000, 32'h4a0},{32'h4000, 32'h4702f000, 32'hbd0},{32'h28d00000, 32'h1081a204, 32'h1278},{32'hc0056000, 32'h34c05420, 32'h140},{32'heaa00000, 32'h1d40e, 32'h3b0},{32'hb8a80000, 32'h3bc00025, 32'h170},{32'hd0020000, 32'h8b000002, 32'ha60},{32'h16720402, 32'h52c0000e, 32'he98},{32'h40000000, 32'h22429414, 32'ha50},{32'he5600000, 32'h33019c0c, 32'h7b8},{32'h8e80000, 32'hae09, 32'h10c0},{32'ha5400080, 32'h2540b01d, 32'h290},{32'haa00000, 32'h5e82381a, 32'h0},{32'h3b180002, 32'h67c00004, 32'hbd8},{32'h80000000, 32'h7f808402, 32'h210},{32'h4e0a000, 32'h1e800000, 32'h12b0},{32'h44c00400, 32'h1580ac15, 32'h178},{32'hba746402, 32'h52020c1a, 32'ha68},{32'h67300000, 32'h1a80e422, 32'haa8},{32'hae00000, 32'h22000000, 32'h440},{32'h34000, 32'h29600, 32'h680},{32'hf0020000, 32'hc, 32'h4a0},{32'h4000, 32'h11840800, 32'h230},{32'h5180000, 32'hb212, 32'hbd0},{32'h45400000, 32'h12000002, 32'h260},{32'h7500090, 32'h80c05600, 32'h0},{32'h0, 32'h21008600, 32'h760},{32'h4c00410, 32'hae00, 32'hee8},{32'h0, 32'h5282ae00, 32'h0},{32'h20006000, 32'h1c80d407, 32'h0},{32'h7280080, 32'h2240e600, 32'h0},{32'h400, 32'h10808400, 32'h688},{32'he0046010, 32'h79012a02, 32'h180},{32'had00000, 32'hc808c00, 32'h220},{32'h4e00000, 32'h11c42000, 32'h0},{32'h1300000, 32'h5ec1c400, 32'h5a0},{32'h8b00000, 32'h52829400, 32'h268},{32'h46000, 32'h2201d800, 32'h460},{32'hc8800030, 32'h1c039e06, 32'h380},{32'hb5580402, 32'h14, 32'hd58},{32'h0, 32'he400, 32'h12d0},{32'h8800000, 32'h0, 32'ha90},{32'h24700410, 32'h11808604, 32'h1268},{32'h7700000, 32'h6020, 32'h140},{32'h5aa00000, 32'h20, 32'h188},{32'h20000000, 32'h29008e0a, 32'h1080},{32'h4a980000, 32'h15, 32'hbe8},{32'h3a700010, 32'h8482960e, 32'h510},{32'h6b00000, 32'h3b039c00, 32'h0},{32'h7000000, 32'h9381a400, 32'h690},{32'hc4e00000, 32'h1c41dc0e, 32'h470},{32'haaa00000, 32'h1c800006, 32'h3a0},{32'h37500000, 32'h3c845207, 32'h6f0},{32'hd6b00000, 32'h54c2941a, 32'h0},{32'hd0000008, 32'h1d, 32'h248},{32'h60000000, 32'h3a806225, 32'h740},{32'h5580000, 32'ha, 32'h520},{32'h5400000, 32'h1600b000, 32'hee0},{32'h96a00000, 32'h24, 32'hab8},{32'h50000000, 32'h2380000a, 32'h1150},{32'h4c00000, 32'h34800000, 32'h680},{32'h86800000, 32'h25, 32'h770},{32'h65400000, 32'h11008c03, 32'h0},{32'h67600000, 32'h1400a805, 32'h3a8},{32'h38e80000, 32'h3a01200f, 32'h750},{32'h7100000, 32'h2d83f000, 32'h5c0},{32'h7100000, 32'h9, 32'heb0},{32'h45400000, 32'h3981c80a, 32'h6e0},{32'ha89d0000, 32'h29429c14, 32'h2d0},{32'h49720000, 32'hc00b220, 32'h170},{32'ha980000, 32'h1c04ac07, 32'h770},{32'h5056000, 32'h3b011000, 32'h780},{32'ha7100000, 32'h2501a625, 32'h0},{32'hcac00000, 32'h24, 32'hf40},{32'h4a800000, 32'h1580b424, 32'h2e0},{32'h9506000, 32'h2501d000, 32'h0},{32'h8c00000, 32'h2c816c00, 32'h0},{32'h8c00000, 32'h12800, 32'h12c0},{32'h55000402, 32'h2901480a, 32'h1238},{32'h46410, 32'h39c3a200, 32'h2d8},{32'h0, 32'h45003, 32'ha88},{32'h18750002, 32'hc417007, 32'h1230},{32'hf8b00000, 32'h3d839c0e, 32'h7b0},{32'he5180000, 32'h3b81280e, 32'h788},{32'h47280000, 32'hf81de04, 32'h0},{32'h7ac00402, 32'h5, 32'hfc8},{32'ha0000000, 32'h8980e006, 32'h2e8},{32'h67600000, 32'h7e80000b, 32'h758},{32'hac00000, 32'h0, 32'h1270},{32'h4700010, 32'h3ac14a00, 32'h0},{32'h40000000, 32'h1a40a, 32'h1270},{32'h15600002, 32'h2001ec03, 32'h11b0},{32'he4e00000, 32'h1d429414, 32'h1030},{32'hb5280000, 32'h700380b, 32'h11a0},{32'hc6a00000, 32'h3dc2e40b, 32'hba0},{32'hf9500000, 32'h7f80000e, 32'h230},{32'h44c00000, 32'h3980000e, 32'h6f0},{32'haa980000, 32'h1b000006, 32'h370},{32'h7500000, 32'h2e00e200, 32'h0},{32'he0030000, 32'h80806002, 32'h5c8},{32'h1ae00000, 32'h7501cc0d, 32'h730},{32'h24e00000, 32'h3880000d, 32'h730},{32'h44f50000, 32'h1a60f, 32'hf70},{32'h8a800000, 32'h79000004, 32'h250},{32'hfad00000, 32'h67800014, 32'h910},{32'he6b00000, 32'h73803a0b, 32'h10e8},{32'h7400000, 32'h11800000, 32'h1260},{32'h6800000, 32'he, 32'h730},{32'h5400000, 32'hd823, 32'h0},{32'ha708090, 32'h2e449200, 32'h0},{32'h40000000, 32'hb800002, 32'h160},{32'h25580000, 32'h17006205, 32'h1000},{32'h35580002, 32'h5701ce0d, 32'hd50},{32'h76b00000, 32'h8d80000e, 32'h7b0},{32'h24c00000, 32'h3d40d, 32'h750},{32'hf9500000, 32'h1d, 32'h258},{32'h0, 32'h6882f600, 32'h0},{32'h60f00000, 32'h4, 32'hba8},{32'h80050000, 32'h16008e05, 32'hfc0},{32'h6a80400, 32'h39c00000, 32'h378},{32'h20000000, 32'h3984900e, 32'h5e8},{32'h4b180000, 32'h2e805423, 32'h5e0},{32'hab026000, 32'h2e80ac0b, 32'h2e0},{32'h45056000, 32'he022, 32'h370},{32'hdaa00100, 32'h8a408c15, 32'h240},{32'h28000, 32'h3a81ee00, 32'h0},{32'h40030000, 32'h5b02d41e, 32'h758},{32'h9580000, 32'h54800000, 32'h0},{32'h76700002, 32'h2ea04, 32'h0},{32'he0000000, 32'h1280b01d, 32'h170},{32'h2a988000, 32'h1e40f, 32'he90},{32'he8a80000, 32'h5c01cc16, 32'h310},{32'ha9c0400, 32'h39c00000, 32'h5e8},{32'hb0000002, 32'hbc0000b, 32'h2d0},{32'ha0b00000, 32'h17400004, 32'h0},{32'h6a700400, 32'h3980e20e, 32'h248},{32'he0056080, 32'h3ac04001, 32'h1090},{32'hcaa00000, 32'hb806c02, 32'hb60},{32'he503a000, 32'h3a81dc0e, 32'h0},{32'h8e80000, 32'h3c02a600, 32'h0},{32'h96700002, 32'h5e82f405, 32'hd00},{32'h6a00000, 32'h12c00000, 32'hf28},{32'h30000010, 32'h1ce0f, 32'h0},{32'h20000000, 32'h5c440c01, 32'hf0},{32'h29500000, 32'h1c00e00f, 32'h0},{32'hd0046050, 32'h46a05, 32'h0},{32'h70000002, 32'h1340000e, 32'h0},{32'h60000000, 32'h1, 32'h100},{32'h45400080, 32'hbc3ac17, 32'hba0},{32'hf5280000, 32'h5b43721b, 32'h780},{32'hf0020000, 32'hb80600e, 32'h180},{32'h24e00000, 32'h5c01e21a, 32'h320},{32'haa980000, 32'h4882f617, 32'hbd0},{32'h64e80000, 32'h1801024, 32'h0},{32'hae00000, 32'hf, 32'h0},{32'ha700010, 32'he200, 32'hf8},{32'hc0000000, 32'h7049c01, 32'h0},{32'h7280000, 32'h8002c00, 32'h100},{32'h5180000, 32'h5d02e400, 32'h5f0},{32'h8980000, 32'h13004203, 32'hf20},{32'h55580400, 32'he837017, 32'h788},{32'ha8f00000, 32'hc00241e, 32'hb50},{32'heb106000, 32'h1882e016, 32'h0},{32'h2ae00000, 32'h5c401400, 32'h70},{32'hb9500000, 32'h2800017, 32'h0},{32'h60030000, 32'h7001220, 32'hf0},{32'h7500000, 32'h3a600, 32'h798},{32'h0, 32'h3800, 32'hd0},{32'h8800000, 32'h85000002, 32'h10a0},{32'h74e80000, 32'h8434421, 32'hba0},{32'h5000000, 32'h3d81ec00, 32'h780},{32'h6a00000, 32'h13401000, 32'h50},{32'hd0028410, 32'h6216, 32'hf38},{32'ha0000000, 32'h5e833c17, 32'hb58},{32'he7280000, 32'h7c82e200, 32'h90},{32'had00090, 32'h2c3f600, 32'h78},{32'h0, 32'h6803800, 32'h0},{32'h8c00000, 32'h8a00e400, 32'h3a0},{32'h8d00000, 32'h6003400, 32'hf50},{32'hd4e00000, 32'h42801, 32'hc0},{32'h8800000, 32'h18c00, 32'h0},{32'h61300000, 32'h5d43b20f, 32'h0},{32'h50400, 32'h1ee00, 32'h58},{32'h0, 32'h7782d800, 32'hef0},{32'h4e00000, 32'h2f400, 32'h940},{32'h8800000, 32'h1400b824, 32'h0},{32'h6ae00000, 32'h3d04680e, 32'h98},{32'hc9580000, 32'h7c009001, 32'h260},{32'h28d0a000, 32'he007, 32'h0},{32'h8b000000, 32'h3c03a001, 32'h7a0},{32'h710a000, 32'h8000000, 32'hd60},{32'h86800000, 32'h71802c15, 32'h0},{32'h77280002, 32'hf, 32'hbb8},{32'h0, 32'h2a415, 32'hf30},{32'h6aa00000, 32'h5b00000f, 32'h1d0},{32'h6801400, 32'h25800, 32'hcc8},{32'hb1300000, 32'h5501cc17, 32'haa0},{32'he5180000, 32'h5300ba14, 32'hcc0},{32'h86a80400, 32'h3d405404, 32'hf8},{32'hab000000, 32'h1d00b805, 32'h2a0},{32'haa30090, 32'h87403600, 32'h3a8},{32'h0, 32'h55835803, 32'h7a8},{32'h19580000, 32'h56002802, 32'had0},{32'h97100000, 32'h3037815, 32'h60},{32'h5180000, 32'h74800007, 32'h7a0},{32'hc7500000, 32'h2a61e, 32'h0},{32'he1700000, 32'h182da00, 32'h80},{32'hcad00000, 32'h5f42d816, 32'hdd0},{32'hf8a80000, 32'h5540001a, 32'ha80},{32'hf0020000, 32'h54029c14, 32'ha60},{32'h8980080, 32'h1d400000, 32'h268},{32'he0000000, 32'hb80ba1d, 32'h260},{32'h2ad00000, 32'h4, 32'ha90},{32'h65400000, 32'h2b001, 32'h0},{32'h49400000, 32'h80181f, 32'h0},{32'hae00000, 32'h3400000, 32'hfd8},{32'h80000000, 32'h2000c00, 32'h7a8},{32'hc7280000, 32'h4001c21, 32'hb78},{32'h39580000, 32'h1f, 32'h88},{32'hd0000410, 32'h32e16, 32'ha88},{32'he0000000, 32'h1d03a414, 32'h7a0},{32'h68d0a000, 32'hb805, 32'h2e0},{32'h5600000, 32'h12806000, 32'h0},{32'hc7000000, 32'h1a, 32'h240},{32'h8a800000, 32'h3dc15, 32'h0},{32'hab000000, 32'h1000000, 32'h0},{32'hcac00000, 32'h5702b81d, 32'h0},{32'h7600000, 32'h5c001000, 32'hd10},{32'he6b08000, 32'hc00, 32'h0},{32'hb000000, 32'h5c02e000, 32'he50},{32'h6a00000, 32'h8004000, 32'hd0},{32'h6a00090, 32'h5443ba00, 32'h0},{32'h80000000, 32'h17000005, 32'h7a8},{32'h7400000, 32'h641f, 32'h0},{32'h6b000000, 32'he, 32'haa0},{32'h5400000, 32'h7501e400, 32'h7a0},{32'h98d00000, 32'h1a, 32'had8},{32'hc0000000, 32'h10001a16, 32'hb70},{32'h9ad00002, 32'h2ba00, 32'hd48},{32'h10000000, 32'h4a02f417, 32'hbe0},{32'ha8d00000, 32'h4400006, 32'h0},{32'h51700000, 32'h2e21c, 32'h0},{32'h90000000, 32'h4221, 32'h0},{32'hc0000000, 32'h5d02e805, 32'h630},{32'h86a50000, 32'h400ba00, 32'h80},{32'h45580000, 32'h3183b017, 32'h268},{32'h28e80000, 32'h55c1cc0f, 32'h0},{32'h6b000000, 32'h3e004, 32'h260},{32'h29500000, 32'h4, 32'h0},{32'h1700000, 32'h1a82e017, 32'hb78},{32'ha8e80000, 32'h4b01ec17, 32'h7c0},{32'hac28000, 32'h55820c00, 32'hd80},{32'h65180000, 32'h5cc0181a, 32'h60},{32'h5600000, 32'h3c800, 32'h0},{32'hd8700002, 32'h86803c05, 32'hb0},{32'h6a00000, 32'h7642ea00, 32'h0},{32'h0, 32'h443ea00, 32'h0},{32'h50000000, 32'h5402ac17, 32'hab0},{32'h4e00000, 32'h13000000, 32'h7a8},{32'h40030000, 32'h76019017, 32'h268},{32'he7280000, 32'h5fc31418, 32'h0},{32'h18680400, 32'h38e17, 32'h7c8},{32'hc0000000, 32'h7d001400, 32'hbe8},{32'hc8e80000, 32'h55c1e005, 32'h7a0},{32'h49500000, 32'h55801a15, 32'hd50},{32'hca980000, 32'h1842b815, 32'ha80},{32'he8a80000, 32'h5f003e12, 32'hbe0},{32'h5580000, 32'h87003c00, 32'h10e0},{32'h84e00000, 32'h3001800, 32'h0},{32'hd7600082, 32'h1342ae19, 32'h0},{32'h0, 32'h19800, 32'h0},{32'h51300000, 32'h32817, 32'hff0},{32'h5000000, 32'h53000000, 32'h7c0},{32'h6b00000, 32'h69800000, 32'h60},{32'h4c00000, 32'h3d004002, 32'hf0},{32'hc8ab0000, 32'h2a419, 32'h7a8},{32'h9400000, 32'h8842c00, 32'h100},{32'hd5180000, 32'h58037815, 32'hb00},{32'hf5180000, 32'h5f431419, 32'hcc0},{32'he8b00000, 32'h4c803e19, 32'h0},{32'haf00000, 32'h5c801a17, 32'h370},{32'hca980000, 32'h3c01, 32'h0},{32'h4a000, 32'h5dc3f800, 32'hc20},{32'he8800000, 32'h5682b014, 32'hc0},{32'h898a000, 32'h3000000, 32'h50},{32'h6800090, 32'h3d433a00, 32'h0},{32'h10000000, 32'h602b002, 32'haf0},{32'h68d00000, 32'h55c03421, 32'h0},{32'heb000000, 32'h102c015, 32'h0},{32'hae00000, 32'h58432c00, 32'h0},{32'hb1300000, 32'h1800bc18, 32'hfe8},{32'h38000, 32'h70c2fa00, 32'h0},{32'h10, 32'h5cc03e00, 32'h0},{32'h80000000, 32'h3c24, 32'h0},{32'hfa700210, 32'h7042a218, 32'h0},{32'h0, 32'h56c01800, 32'h0},{32'he0008000, 32'h5583381a, 32'h0},{32'h8b180000, 32'h3415, 32'h0},{32'h8b000000, 32'h3c21, 32'h0},{32'h6b000000, 32'h2a01a, 32'hb00},{32'ha5400200, 32'h6a43b818, 32'h0},{32'h4b300080, 32'h1842f814, 32'hc68},{32'h9700000, 32'h70828800, 32'hc60},{32'h87300100, 32'h7f42e80c, 32'hbb0},{32'h89500000, 32'h56800015, 32'hd60},{32'hea980000, 32'h5b80741b, 32'hac8},{32'hdb180402, 32'h0, 32'hd38},{32'h0, 32'h32c00, 32'hab0},{32'h85000000, 32'h3c1a, 32'h0},{32'hb000000, 32'h5c038802, 32'hb90},{32'h8710a000, 32'h58000000, 32'h0},{32'h87400000, 32'h62031019, 32'h0},{32'h87600000, 32'h63402816, 32'hb50},{32'hab100000, 32'h3833400, 32'hbf8},{32'hdb180000, 32'h17, 32'hcf8},{32'h20000000, 32'h5a82d001, 32'hbb8},{32'h9580000, 32'h56c2d800, 32'he00},{32'h88800000, 32'h5680001a, 32'hf0},{32'h4a980000, 32'h3302ac17, 32'hbb0},{32'haad40000, 32'h55c26415, 32'h0},{32'h4b000080, 32'h8c0d41c, 32'h0},{32'hb000000, 32'h69800016, 32'hb00},{32'h4e80000, 32'h5582c200, 32'hac0},{32'hf0026000, 32'h6a031222, 32'hd40},{32'h14f00000, 32'h21, 32'hb58},{32'hc0000000, 32'h3c29417, 32'hbf0},{32'hb100000, 32'h21, 32'hf0},{32'hca800000, 32'h8016, 32'h0},{32'h6b000000, 32'h55800015, 32'h0},{32'h50056012, 32'h56c2ae1a, 32'h0},{32'h90000000, 32'h6a83541d, 32'hbb8},{32'hc7000000, 32'h56838c06, 32'h0},{32'h9400030, 32'h58035200, 32'h50},{32'hb6800402, 32'h1c, 32'hac8},{32'hc0000000, 32'h15, 32'hac0},{32'h8a800000, 32'h5d80001d, 32'h680},{32'h8a980000, 32'h380001f, 32'h40},{32'h4a980000, 32'h5880001a, 32'hbf8},{32'h7700000, 32'h5ac00000, 32'he18},{32'h70000402, 32'h5bc00015, 32'hce8},{32'h0, 32'h5b808400, 32'hb70},{32'h5180000, 32'h8835000, 32'h0},{32'hc8c00000, 32'h15, 32'hce0},{32'hab00000, 32'h68400000, 32'hb98},{32'h10000000, 32'h7d002016, 32'hfa0},{32'h4e00000, 32'h5c80e000, 32'hb90},{32'h25180000, 32'h2be0d, 32'h0},{32'h1700000, 32'h5dc3f400, 32'hfd0},{32'h25000000, 32'h33416, 32'h10f0},{32'hd5280000, 32'h2c61c, 32'h0},{32'h0, 32'h63830400, 32'hc70},{32'h65180000, 32'h4, 32'h0},{32'hb1700000, 32'h5bc00019, 32'h0},{32'h0, 32'h68000007, 32'haf8},{32'h7700000, 32'h57c2c016, 32'hd30},{32'he8a80000, 32'h69800000, 32'h0},{32'haac00000, 32'h5700001a, 32'haf0},{32'h67500000, 32'h5cc34215, 32'hc60},{32'ha5700000, 32'h5f82ee19, 32'h240},{32'haa980000, 32'h3c00800, 32'h70},{32'h3b100000, 32'h3a82ec16, 32'h0},{32'h28f00000, 32'h31c18, 32'hc70},{32'h5600000, 32'h63c3fe00, 32'h0},{32'h80000000, 32'h6202de18, 32'h1060},{32'h6a80000, 32'h1d034000, 32'h0},{32'h8c00000, 32'h3801800, 32'h0},{32'h10038000, 32'h34a16, 32'h0},{32'h20000000, 32'h280221f, 32'h90},{32'haad00000, 32'h5880001c, 32'haf8},{32'ha7700000, 32'h7831a01, 32'ha0},{32'ha980000, 32'h5fc01800, 32'h0},{32'h8000, 32'h0, 32'h780},{32'h70b00000, 32'h63800017, 32'hc30},{32'h6800000, 32'h5402b800, 32'haf0},{32'h8d00000, 32'h31000, 32'hc30},{32'h28800000, 32'h201f, 32'h50},{32'haa00080, 32'h3c00000, 32'hbc8},{32'hc0000000, 32'h5f82dc19, 32'h0},{32'h9580000, 32'h383e800, 32'h0},{32'h8c00000, 32'h82cc00, 32'hb40},{32'hc8d00000, 32'h62845c22, 32'hb28},{32'hb180400, 32'h7c00000, 32'h78},{32'h0, 32'h61030c00, 32'hcd0},{32'hc4e00000, 32'h5e433018, 32'hc80},{32'h6b100000, 32'h5e031e0f, 32'hbf0},{32'h47500000, 32'h64032419, 32'haf8},{32'h97600000, 32'h64830418, 32'hc90},{32'h45180000, 32'h7802201, 32'he0},{32'h5580000, 32'h33800, 32'hbc0},{32'hc5000000, 32'h2ac15, 32'haf0},{32'h6b100000, 32'h1000016, 32'h98},{32'hcac00000, 32'h4002000, 32'h0},{32'he7600000, 32'h62c2a018, 32'hfe0},{32'h45280000, 32'h6302ac18, 32'hc60},{32'h518a000, 32'h6103f800, 32'h70},{32'h8c00100, 32'h69401c01, 32'hec0},{32'h28a80000, 32'h65032819, 32'hbf8},{32'h7280000, 32'h64032600, 32'hca0},{32'hc7500000, 32'h64c00001, 32'hcb8},{32'ha000a000, 32'h14, 32'hcf0},{32'h25400000, 32'h7c82bc16, 32'hb00},{32'h44ec0000, 32'h59830019, 32'haf8},{32'he7600000, 32'h3201f, 32'hb48},{32'hae00000, 32'h7f002200, 32'hac0},{32'h6800010, 32'h57830e00, 32'haf0},{32'hf0034000, 32'h63402024, 32'h90},{32'he0028000, 32'h62830c22, 32'hc88},{32'h1b180000, 32'h65800001, 32'hc20},{32'he6800000, 32'h86000001, 32'h110},{32'had00080, 32'h7c00000, 32'hca8},{32'h0, 32'h32c00, 32'hbf0},{32'hc5000010, 32'h5a02be00, 32'hb40},{32'h35580000, 32'h60000016, 32'h0},{32'h20006000, 32'h5803f416, 32'h0},{32'h7280000, 32'h4032201, 32'h70},{32'hf6a80080, 32'h57c00018, 32'h0},{32'he0000400, 32'h57831824, 32'h98},{32'h8ae00000, 32'h61831018, 32'hc50},{32'h8d0a000, 32'h61800000, 32'hcb0},{32'h4c00000, 32'h7804000, 32'h0},{32'h8c00000, 32'h7002fc00, 32'hb50},{32'hc4e00000, 32'h2bc1c, 32'hb20},{32'h2b100000, 32'h5fc32418, 32'hc90},{32'h5600010, 32'h5a430200, 32'h0},{32'h0, 32'h382c000, 32'h0},{32'he8c00000, 32'h6302bc18, 32'h0},{32'h17280000, 32'h63830c01, 32'hc80},{32'h7100000, 32'h2001, 32'h0},{32'h80058080, 32'h62c31a18, 32'h0},{32'he000a000, 32'h3800017, 32'hb40},{32'h34e80000, 32'h782b419, 32'had0},{32'h4e00000, 32'h0, 32'h118},{32'h0, 32'h2fe02, 32'h110},{32'h2a000, 32'h0, 32'hb28},{32'h0, 32'h5e032618, 32'h7c0},{32'h6a80000, 32'h34800, 32'h90},{32'h8800000, 32'h6183fc00, 32'h0},{32'h8c00000, 32'h62831c00, 32'h0},{32'h18c00012, 32'h45a01, 32'h0},{32'h400, 32'h0, 32'hc58},{32'h0, 32'h5a000000, 32'h90},{32'h6800000, 32'h882fc00, 32'he10},{32'h4e00000, 32'h5982b600, 32'hc10},{32'h7500400, 32'h0, 32'h118},{32'h0, 32'h64832400, 32'hc30},{32'h6a00000, 32'h2a000, 32'hbf0},{32'h5000000, 32'h58800000, 32'hce0},{32'h6800000, 32'h31c00, 32'hc50},{32'ha8800000, 32'h2cc16, 32'hec0},{32'h8a80000, 32'h0, 32'hc88},{32'h0, 32'h33019, 32'hca0},{32'hb100000, 32'h5f800000, 32'hce0},{32'h26800000, 32'h5f00001c, 32'h0},{32'h7400000, 32'h66033000, 32'h0},{32'h7000000, 32'h5682b400, 32'h110},{32'h6a00000, 32'h6902c000, 32'hb10},{32'h8d00000, 32'h5f832600, 32'hac0},{32'h6800000, 32'h5782c400, 32'h0},{32'h28c00000, 32'h32419, 32'hc50},{32'hf8a80000, 32'h66800818, 32'h0},{32'h87000000, 32'h1480b, 32'h1010},{32'h5280000, 32'h61046c00, 32'h0},{32'ha8c00000, 32'h4a003, 32'h1e0},{32'hfb100000, 32'h70800017, 32'ha30},{32'h6800000, 32'h60000000, 32'h0},{32'he0006000, 32'he000020, 32'h1a0},{32'h6a980000, 32'h2b618, 32'hc40},{32'had00000, 32'h0, 32'hb18},{32'h10000000, 32'h18, 32'hb20},{32'h30020000, 32'h16, 32'h0},{32'h30000000, 32'h69000019, 32'hb40},{32'h4c00000, 32'h34801, 32'hb10},{32'h99500000, 32'h64830c0b, 32'h0},{32'h7000000, 32'h0, 32'h0},{32'h0, 32'h0, 32'h1e8},{32'h400, 32'h2fe00, 32'hc18},{32'hc0000000, 32'h2fc17, 32'ha60},{32'haa00000, 32'he400000, 32'h0},{32'h0, 32'h0, 32'hc48},{32'h400, 32'h0, 32'hb28},{32'he0000000, 32'h31818, 32'hb20},{32'h8a80000, 32'h5a045800, 32'h0},{32'h7000000, 32'h0, 32'h0},{32'h0, 32'h62832400, 32'hb18},{32'h8c00000, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h54000000, 32'hbf0},{32'h4c00000, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'hc80},{32'hf0020000, 32'h2d018, 32'ha0},{32'h8800000, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'hca8},{32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h40000000, 32'h5f80001a, 32'h0},{32'h7400000, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h480, 32'h8cc00000, 32'hc88},{32'h0, 32'h8a800000, 32'h1170},{32'h26800000, 32'h8c800019, 32'hca0},{32'had00000, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h2fe00, 32'he68},{32'he0000000, 32'h5782fc17, 32'h0},{32'h8e80000, 32'h2bc18, 32'he60},{32'h5280000, 32'h0, 32'h0},{32'h0, 32'h7800000, 32'hb50},{32'h4c00000, 32'h0, 32'h0},{32'h0, 32'h0, 32'hca8},{32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'hf0000000, 32'h73400017, 32'h0},{32'h10000000, 32'h18, 32'h0},{32'h0, 32'h5a800000, 32'h110},{32'h6800000, 32'h73000018, 32'hb20},{32'h6a80000, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h2d400, 32'h1a0},{32'h8800000, 32'h0, 32'h0},{32'h10000000, 32'h18, 32'h0},{32'h0, 32'h60000018, 32'h0},{32'h56000, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0},{32'hb0000000, 32'h16, 32'h0},{32'h0, 32'h0, 32'h0},{32'h10000002, 32'h18, 32'h0},{32'h0, 32'h0, 32'h0},{32'h1, 32'h0, 32'h0}};

