//Constant array to load the A matrix
localparam integer A_size = 665;
localparam integer A[0:664] = '{32'h3e088c61, 32'hbd8888b5, 32'hb76ae18b, 32'hbd8888b5, 32'h3e088c61, 32'hbd8888b5, 32'hb76ae18b, 32'hbd8888b5, 32'h3e088ace, 32'hbd8888b5, 32'hbd8888b5, 32'hb70637bd, 32'h4170021b, 32'hb9fa9c13, 32'hb58637bd, 32'hb796feb5, 32'hb796feb5, 32'hb9fb224b, 32'h3b272eae, 32'hb8b88ca4, 32'hba828c37, 32'hba81a155, 32'hbd8888b5, 32'hbd8888b5, 32'h360637bd, 32'h390b75ea, 32'h3eaad2fe, 32'hb9712c28, 32'hbe4ccccd, 32'hb95f58c1, 32'hb76ae18b, 32'hb78637bd, 32'hbab02928, 32'h39ad8a11, 32'h3c51dcd7, 32'hbc441dd2, 32'h3955e8d5, 32'h3e08900c, 32'hbd8888b5, 32'hb7f34507, 32'hbd8888b5, 32'h3e088bdb, 32'hbd8888b5, 32'hbd8888b5, 32'hb75a1a93, 32'h40f00560, 32'hba19e0e7, 32'hb58637bd, 32'hb816feb5, 32'hb80a697b, 32'hba1aaa3b, 32'h3b81450f, 32'hba2d46f6, 32'hbad6909b, 32'hba8a8b09, 32'hbd8888b5, 32'hbd8888b5, 32'h368637bd, 32'h3948472c, 32'h3eaae4d2, 32'hb9d23d4f, 32'hbe4ccccd, 32'hb9798fa3, 32'hb7f34507, 32'hb81f6230, 32'hbb6874c9, 32'h3966afcd, 32'h3cd55821, 32'hbcc41dd2, 32'h3aa91538, 32'h3e088c61, 32'hb76ae18b, 32'hbd8888b5, 32'h3e088ace, 32'hbd8888b5, 32'hb716feb5, 32'h3cf3c2db, 32'hb87fda40, 32'hb58637bd, 32'hbcf2c301, 32'hb87fda40, 32'hb76ae18b, 32'hb8a5accd, 32'h3c69680e, 32'h3851b717, 32'hb78e9b39, 32'hbb113a50, 32'hbd8888b5, 32'hbd8888b5, 32'h36c9539c, 32'hb76ae18b, 32'h3eaaad1d, 32'h358637bd, 32'hb749539c, 32'hbcf2c301, 32'hb796feb5, 32'h3f5cedc4, 32'hb796feb5, 32'hbf555550, 32'h3d13165d, 32'hbcc41dd2, 32'hbc441dd2, 32'h3e08900c, 32'hbd8888b5, 32'hbd8888b5, 32'hb7f34507, 32'h3f800000, 32'hbd8888b5, 32'h3e088bdb, 32'hbd8888b5, 32'hb75a1a93, 32'hbd8888b5, 32'hbe4ccccd, 32'hbd8888b5, 32'h3eaaaf14, 32'hb6a7c5ac, 32'hb80a697b, 32'h36a7c5ac, 32'hb7f34507, 32'hbcc41dd2, 32'h358637bd, 32'h3cc4d445, 32'hb58637bd, 32'hb80e9b39, 32'hb7c9539c, 32'hb80637bd, 32'hb79f6230, 32'h3b8c2614, 32'hbb8b08dd, 32'h378e9b39, 32'hb80e9b39, 32'hbb8b08dd, 32'h3ed78983, 32'hb7e27e0f, 32'hbed55561, 32'hbcc41dd2, 32'hb75a1a93, 32'hb60637bd, 32'hb7e27e0f, 32'h3cc475e6, 32'hb716feb5, 32'hb851b717, 32'hbb0e25c8, 32'hb88e9b39, 32'hb7a7c5ac, 32'hbc441dd2, 32'h3c6a0ba2, 32'h3f800000, 32'h3e088c61, 32'hb76ae18b, 32'hbd8888b5, 32'hb76ae18b, 32'h3c449fd8, 32'hb78637bd, 32'h3e088a48, 32'hbd8888b5, 32'hb6c9539c, 32'h3bd6c2f0, 32'hb716feb5, 32'hb727c5ac, 32'hbbd6238e, 32'hbd8888b5, 32'hbd8888b5, 32'hb79f6230, 32'h3eaaad1d, 32'hb6c9539c, 32'hb727c5ac, 32'h3c449ba6, 32'hb76ae18b, 32'hbc441dd2, 32'hbf555550, 32'hb78637bd, 32'hbbd6238e, 32'hb76ae18b, 32'h3f57038e, 32'h40055554, 32'hbf555550, 32'h3f800000, 32'hbed55561, 32'hbf555550, 32'hbd8888b5, 32'h3e08900c, 32'hbd8888b5, 32'hb7f34507, 32'hbd8888b5, 32'h3e088d2a, 32'hbd8888b5, 32'hb796feb5, 32'hbe4ccccd, 32'hbd8888b5, 32'hbd8888b5, 32'h3eaaaf79, 32'hb7da1a93, 32'h377ba882, 32'hb7da1a93, 32'hbcc41dd2, 32'hb7f34507, 32'h38e27e0f, 32'h3ccfd8f1, 32'hb910b418, 32'hbaaf5fd4, 32'hb812ccf7, 32'hb6c9539c, 32'hb8e8c8ac, 32'h3c8f861a, 32'hb8e8c8ac, 32'hbc8da7f4, 32'hb796feb5, 32'hb910b418, 32'hbaa15981, 32'hb8dc3372, 32'h3cd0a244, 32'hb816feb5, 32'hbcc41dd2, 32'hbed55561, 32'hb816feb5, 32'hbc8da7f4, 32'hb816feb5, 32'h3ede392e, 32'h3cc41dd2, 32'hbc441dd2, 32'hbc441dd2, 32'h3e088c61, 32'hb76ae18b, 32'hbd8888b5, 32'hbc441dd2, 32'hb76ae18b, 32'h3c449fd8, 32'hb78637bd, 32'h3e088a48, 32'hb6eae18b, 32'hbd8888b5, 32'h3bd66f0d, 32'hb60637bd, 32'hb78637bd, 32'hbbd5cfab, 32'hb6eae18b, 32'h3c447a18, 32'hb60637bd, 32'hb76ae18b, 32'hbc441dd2, 32'hbd8888b5, 32'hbd8888b5, 32'hb79f6230, 32'h3eaaad1d, 32'hbf555550, 32'hb78637bd, 32'hbbd5cfab, 32'hb76ae18b, 32'h3f5702f7, 32'h3e088c61, 32'hb76ae18b, 32'hbd8888b5, 32'h3e088ace, 32'hbd8888b5, 32'hb716feb5, 32'h3cf02c4d, 32'hb896feb5, 32'hb60637bd, 32'hbceef805, 32'hb8991794, 32'hb76ae18b, 32'hb8dc3372, 32'h3c698138, 32'h385a1a93, 32'hb77ba882, 32'hbb101d19, 32'hbd8888b5, 32'hbd8888b5, 32'h36c9539c, 32'hb77ba882, 32'h3eaaad1d, 32'h3649539c, 32'hb749539c, 32'h3e088c61, 32'hb76ae18b, 32'hbd8888b5, 32'hb76ae18b, 32'h3c449fd8, 32'hb78637bd, 32'h3e088a48, 32'hbd8888b5, 32'hb6c9539c, 32'h3bd6ba8c, 32'hb727c5ac, 32'hb716feb5, 32'hbbd6238e, 32'hbd8888b5, 32'hbd8888b5, 32'hb79f6230, 32'h3eaaad1d, 32'hb6c9539c, 32'hb716feb5, 32'h3c449774, 32'hb76ae18b, 32'hbc441dd2, 32'hb78637bd, 32'hbbd6238e, 32'hb76ae18b, 32'h3f57038e, 32'hbf555550, 32'h3f800000, 32'h3e088c61, 32'hb76ae18b, 32'hbd8888b5, 32'hb76ae18b, 32'h3c449fd8, 32'hb78637bd, 32'h3bd6a9c5, 32'hb79f6230, 32'hbbd60a63, 32'h3e088a48, 32'hbd8888b5, 32'hb6eae18b, 32'hbd8888b5, 32'hb79f6230, 32'hbd8888b5, 32'h3eaaad1d, 32'hb6eae18b, 32'h3c4471b4, 32'hbc441dd2, 32'hb76ae18b, 32'hbc441dd2, 32'h3cc41dd2, 32'hbc441dd2, 32'hbf555550, 32'hb78637bd, 32'hbbd60a63, 32'hb76ae18b, 32'h3f57035c, 32'hbf555550, 32'h40055554, 32'hbf555550, 32'h3f800000, 32'hbed55561, 32'hbd8888b5, 32'h3e08900c, 32'hbd8888b5, 32'hb7f34507, 32'hbd8888b5, 32'h3e088d2a, 32'hbd8888b5, 32'hb796feb5, 32'hbe4ccccd, 32'hbd8888b5, 32'hbd8888b5, 32'h3eaaaf79, 32'hb7f34507, 32'h377ba882, 32'hb7c0f020, 32'hbcc41dd2, 32'hb7f34507, 32'h38e06530, 32'h3ccfce74, 32'hb910b418, 32'hbaae9681, 32'hb812ccf7, 32'hb6c9539c, 32'hb8e6afcd, 32'h3c8f1b26, 32'hb8e8c8ac, 32'hbc8d3cff, 32'hb796feb5, 32'hb910b418, 32'hbaa04d12, 32'hb8da1a93, 32'h3cd08f65, 32'hb816feb5, 32'hbcc41dd2, 32'hbed55561, 32'hb816feb5, 32'hbc8d3cff, 32'hb816feb5, 32'h3ede327f, 32'hbc441dd2, 32'hbcc41dd2, 32'h3f5e86b6, 32'hbf555550, 32'h3e088b54, 32'hbd8888b5, 32'hb7388ca4, 32'h3e088a48, 32'hbd8888b5, 32'hb6eae18b, 32'hbd8888b5, 32'hbd8888b5, 32'h3eaaac11, 32'hb727c5ac, 32'hb727c5ac, 32'h3b73eccc, 32'hbb734507, 32'h358637bd, 32'hb58637bd, 32'hbb734507, 32'h3f564ae0, 32'hb78e9b39, 32'hb78e9b39, 32'hbf555550, 32'hb6eae18b, 32'hb78e9b39, 32'h3c44827b, 32'hbc441dd2, 32'hbc441dd2, 32'hb7388ca4, 32'hb78e9b39, 32'hb58637bd, 32'h3c449774, 32'hbceef805, 32'hb796feb5, 32'hbf555550, 32'h3f5ccf5b, 32'hb796feb5, 32'hbc441dd2, 32'hb716feb5, 32'hb849539c, 32'hbb0dc11e, 32'hb890b418, 32'hb7b88ca4, 32'h3c69fadb, 32'hbc441dd2, 32'hbcc41dd2, 32'hbf555550, 32'h3f5e86b6, 32'hbc441dd2, 32'h3f5b763e, 32'hbf555550, 32'hbc441dd2, 32'h3e088c61, 32'hb76ae18b, 32'hbd8888b5, 32'h3e088ace, 32'hbd8888b5, 32'hb716feb5, 32'h3cf03afb, 32'hb88205ff, 32'hb58637bd, 32'hbcef3d3a, 32'hb8734507, 32'hb76ae18b, 32'hb8a17b0f, 32'h3c689a89, 32'h384d8559, 32'hb78e9b39, 32'hbb0e1501, 32'hbd8888b5, 32'hbd8888b5, 32'h36c9539c, 32'hb80a697b, 32'h3eaaacfb, 32'h358637bd, 32'h36eae18b, 32'hbcef3d3a, 32'hb796feb5, 32'h3f5cd196, 32'hb796feb5, 32'hbf555550, 32'h3d13165d, 32'hbc441dd2, 32'hbcc41dd2, 32'h3e088c61, 32'hbd8888b5, 32'hb76ae18b, 32'h3e088a48, 32'hbd8888b5, 32'hb6c9539c, 32'hbd8888b5, 32'hbd8888b5, 32'h3eaaacfb, 32'hb796feb5, 32'hb76ae18b, 32'h3c44a83b, 32'hb78e9b39, 32'hb60637bd, 32'hb75a1a93, 32'hb58637bd, 32'h3bd7a56e, 32'hbbd70e6f, 32'hb68637bd, 32'hb78e9b39, 32'hbbd70e6f, 32'h3f570564, 32'hb76ae18b, 32'hbf555550, 32'hbc441dd2, 32'hb6c9539c, 32'hb6a7c5ac, 32'hb76ae18b, 32'h3c4486ad, 32'hbd8888b5, 32'h3e08900c, 32'hbd8888b5, 32'hb7f34507, 32'hbd8888b5, 32'h3e088d2a, 32'hbd8888b5, 32'hb796feb5, 32'hbe4ccccd, 32'hbd8888b5, 32'hbd8888b5, 32'h3eaaaf79, 32'hb7da1a93, 32'h377ba882, 32'hb7da1a93, 32'hbcc41dd2, 32'hb7f34507, 32'h38dc3372, 32'h3ccfe154, 32'hb90d8ec9, 32'hbaafe60c, 32'hb816feb5, 32'hb68637bd, 32'hb8e8c8ac, 32'h3c90752e, 32'hb8e8c8ac, 32'hbc8e9d52, 32'hbcc41dd2, 32'hb796feb5, 32'hb910b418, 32'hbaa1dfb9, 32'hb8dc3372, 32'h3cd0a88f, 32'hb816feb5, 32'hb816feb5, 32'hbc8e9d52, 32'hb816feb5, 32'h3ede4884, 32'hbed55561, 32'hbf555550, 32'hbed55561, 32'h3fa4a287, 32'hbc441dd2, 32'hbcc41dd2, 32'h3cc41dd2, 32'hbc441dd2, 32'hbc441dd2, 32'h3e088c61, 32'hbd8888b5, 32'hb76ae18b, 32'h3e088ace, 32'hbd8888b5, 32'hb716feb5, 32'h3ced373b, 32'hb58637bd, 32'hb8841ede, 32'hb87fda40, 32'hbcec3116, 32'hbd8888b5, 32'hbd8888b5, 32'h36c9539c, 32'h3eaaacfb, 32'hb80205ff, 32'h36a7c5ac, 32'h358637bd, 32'hbc441dd2, 32'hb76ae18b, 32'hb8a9de8b, 32'h384d8559, 32'h3c684ad8, 32'hbb0ca3e8, 32'hb78e9b39, 32'hbc441dd2, 32'hb716feb5, 32'hb855e8d5, 32'hb88a697b, 32'hbb08722a, 32'h3c689eba, 32'hb7a7c5ac, 32'hb716feb5, 32'hb851b717, 32'hbb09a027, 32'hb88a697b, 32'hb7a7c5ac, 32'hbc441dd2, 32'h3c68ea3a, 32'hbf555550, 32'hbcec3116, 32'hb796feb5, 32'hb796feb5, 32'h3f5cb934, 32'hbf555550, 32'hbed55561, 32'hbc441dd2, 32'hbf555550, 32'h4006df33, 32'hbc441dd2, 32'hb75a1a93, 32'hb80a697b, 32'hb649539c, 32'hb58637bd, 32'hb58637bd, 32'hbcc41dd2, 32'h3cc486ad, 32'hb70637bd, 32'hb7b88ca4, 32'hba61f7d7, 32'hba102de0, 32'h39dbad3a, 32'hbc441dd2, 32'h3c54e4c9, 32'hbd8888b5, 32'h3e088ace, 32'hb716feb5, 32'hbd8888b5, 32'hbd8888b5, 32'hbd8888b5, 32'hbd8888b5, 32'hbe4ccccd, 32'hbc441dd2, 32'hbd8888b5, 32'hbd8888b5, 32'hbe4ccccd, 32'hbcc41dd2, 32'hbd8888b5, 32'h401e86b6, 32'hbd8888b5, 32'hbe4ccccd, 32'hbcc41dd2, 32'hbd8888b5, 32'hbd8888b5, 32'hbe4ccccd, 32'hbcc41dd2, 32'hbd8888b5, 32'hbd8888b5, 32'hbe4ccccd, 32'hbcc41dd2, 32'hbd8888b5, 32'hbd8888b5, 32'hbe4ccccd, 32'hbcc41dd2, 32'hbd8888b5, 32'h3f800000, 32'hbc441dd2, 32'hbe4ccccd, 32'h4170022d, 32'hba017fc7, 32'hb796feb5, 32'hb796feb5, 32'hb58637bd, 32'hba01c2e3, 32'h3b28e2e3, 32'hba8333fd, 32'hba82adc5, 32'hb8ae1049, 32'hb76ae18b, 32'hbc441dd2, 32'hb78637bd, 32'hbaac3a86, 32'h3c518d26, 32'h393fe3b0, 32'h39b2c83f, 32'hbc441dd2, 32'hb716feb5, 32'hb7b88ca4, 32'hba6cb74e, 32'h39ea5b53, 32'h3c558c8f, 32'hba1741d1, 32'hbd8888b5, 32'hbe4ccccd, 32'hbd8888b5, 32'h360637bd, 32'h390d8ec9, 32'hb9755de6, 32'hb969d51b, 32'h3eaad491};
localparam integer A_BRAMInd[0:664] = '{0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 0, 1, 2, 3, 4, 5, 7, 8, 9, 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 0, 1, 2, 3, 4, 5, 6, 7, 8, 1, 2, 5, 6, 7, 8, 9, 0, 2, 4, 5, 6, 7, 8, 9, 1, 2, 3, 4, 5, 6, 7, 8, 9, 1, 2, 3, 6, 7, 8, 9, 0, 1, 2, 3, 5, 6, 8, 9, 0, 1, 2, 4, 5, 6, 7, 8, 9, 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 0, 1, 2, 4, 5, 6, 7, 8, 9, 0, 1, 2, 4, 6, 7, 8, 9, 0, 1, 2, 3, 4, 5, 6, 7, 8, 0, 1, 3, 7, 8, 9, 0, 2, 5, 6, 7, 8, 9, 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 0, 1, 2, 3, 5, 6, 7, 8, 9, 0, 1, 2, 3, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 8, 9, 0, 2, 3, 4, 5, 6, 7, 9, 0, 1, 2, 3, 4, 5, 6, 8, 9, 0, 3, 5, 6, 7, 8, 9, 1, 2, 3, 4, 6, 8, 0, 1, 2, 3, 4, 7, 8, 9, 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 0, 1, 2, 3, 4, 5, 7, 0, 2, 3, 4, 5, 6, 7, 8, 9, 0, 1, 2, 3, 6, 7, 8, 9, 0, 1, 2, 3, 4, 5, 6, 9, 0, 3, 4, 6, 9, 0, 1, 4, 5, 7, 8, 9, 0, 4, 5, 6, 7, 8, 9, 1, 3, 5, 8, 0, 4, 5, 6, 7, 8, 9, 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 0, 1, 2, 4, 5, 6, 7, 8, 9, 0, 1, 2, 3, 4, 5, 6, 7, 8, 0, 2, 4, 6, 7, 8, 9, 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 0, 3, 4, 7, 8, 9, 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 0, 1, 2, 3, 4, 6, 7, 8, 9, 0, 1, 3, 4, 5, 6, 7, 8, 1, 2, 3, 4, 5, 6, 7, 8, 9, 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 0, 1, 3, 4, 5, 6, 7, 8, 9, 1, 3, 4, 5, 6, 7, 8, 1, 5, 6, 8, 9, 1, 5, 6, 9, 2, 5, 7, 9, 0, 1, 2, 3, 5, 0, 3, 4, 5, 6, 7, 9, 1, 3, 4, 5, 6, 7, 8, 9, 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 0, 5, 6, 7, 8, 2, 3, 4, 5, 4, 5, 6, 7, 8, 9, 0, 2, 3, 4, 5, 6, 7, 8, 9, 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 0, 5, 6, 7, 8, 9, 0, 1, 2, 3, 4, 5, 6, 7, 8};
localparam integer A_BRAMAddr[0:664] = '{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 13, 13, 13, 13, 13, 13, 13, 13, 13, 14, 14, 14, 14, 14, 14, 14, 15, 15, 15, 15, 15, 15, 15, 15, 16, 16, 16, 16, 16, 16, 16, 16, 16, 17, 17, 17, 17, 17, 17, 17, 18, 18, 18, 18, 18, 18, 18, 18, 19, 19, 19, 19, 19, 19, 19, 19, 19, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 23, 23, 23, 23, 23, 23, 23, 23, 23, 24, 24, 24, 24, 24, 24, 24, 24, 25, 25, 25, 25, 25, 25, 25, 25, 25, 26, 26, 26, 26, 26, 26, 27, 27, 27, 27, 27, 27, 27, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 30, 30, 30, 30, 30, 30, 30, 30, 30, 31, 31, 31, 31, 31, 31, 31, 32, 32, 32, 32, 32, 32, 32, 32, 32, 33, 33, 33, 33, 33, 33, 33, 33, 34, 34, 34, 34, 34, 34, 34, 34, 34, 35, 35, 35, 35, 35, 35, 35, 36, 36, 36, 36, 36, 36, 37, 37, 37, 37, 37, 37, 37, 37, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 41, 41, 41, 41, 41, 41, 41, 42, 42, 42, 42, 42, 42, 42, 42, 42, 43, 43, 43, 43, 43, 43, 43, 43, 44, 44, 44, 44, 44, 44, 44, 44, 45, 45, 45, 45, 45, 46, 46, 46, 46, 46, 46, 46, 47, 47, 47, 47, 47, 47, 47, 48, 48, 48, 48, 49, 49, 49, 49, 49, 49, 49, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 51, 51, 51, 51, 51, 51, 51, 51, 51, 51, 52, 52, 52, 52, 52, 52, 52, 52, 52, 53, 53, 53, 53, 53, 53, 53, 53, 53, 54, 54, 54, 54, 54, 54, 54, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 56, 56, 56, 56, 56, 56, 57, 57, 57, 57, 57, 57, 57, 57, 57, 57, 58, 58, 58, 58, 58, 58, 58, 58, 58, 58, 59, 59, 59, 59, 59, 59, 59, 59, 59, 60, 60, 60, 60, 60, 60, 60, 60, 61, 61, 61, 61, 61, 61, 61, 61, 61, 62, 62, 62, 62, 62, 62, 62, 62, 62, 62, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 64, 64, 64, 64, 64, 64, 64, 64, 64, 65, 65, 65, 65, 65, 65, 65, 66, 66, 66, 66, 66, 67, 67, 67, 67, 68, 68, 68, 68, 69, 69, 69, 69, 69, 70, 70, 70, 70, 70, 70, 70, 71, 71, 71, 71, 71, 71, 71, 71, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 73, 73, 73, 73, 73, 74, 74, 74, 74, 75, 75, 75, 75, 76, 76, 77, 77, 77, 77, 77, 77, 77, 77, 77, 78, 78, 78, 78, 78, 78, 78, 78, 78, 78, 79, 79, 79, 79, 79, 79, 80, 80, 80, 80, 80, 80, 80, 80, 80};

//Constant array to load the instruction BRAM
localparam integer total_instructions = 406;
localparam integer sub_instructions = 14;
localparam integer Inst[0:405][0:13] = '{{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h7000000, 32'h1c000, 32'h0, 32'h0, 32'h6a0001a8, 32'h1a8000, 32'ha80006a0, 32'h1},{32'h0, 32'h0, 32'h0, 32'h11072900, 32'h1ac3, 32'h0, 32'h0, 32'h1c000, 32'h0, 32'h6a000, 32'h720d41c8, 32'h1c8000, 32'hc8000000, 32'h1},{32'h0, 32'h0, 32'h0, 32'h9e8c3980, 32'h1064, 32'h0, 32'h4a00000, 32'h12834, 32'h68, 32'h7c000, 32'h4c0001f0, 32'h130000, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'ha0e66b00, 32'h19b4, 32'h0, 32'h7a00000, 32'h1e825, 32'h0, 32'h14000, 32'h140c8190, 32'h0, 32'h30000000, 32'h1},{32'h0, 32'h0, 32'h0, 32'h33ac49c0, 32'h107a, 32'h0, 32'h6800000, 32'hd015000, 32'h54, 32'h54000, 32'h150, 32'h1f0000, 32'h7c0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h152862c0, 32'h1abb, 32'h0, 32'h1400000, 32'h5c18817, 32'h1f000062, 32'h0, 32'h1f0, 32'h0, 32'h58000000, 32'h0},{32'h0, 32'h0, 32'h0, 32'h2c8d5200, 32'h19be, 32'h0, 32'h0, 32'h1e800, 32'h5018030, 32'h64000, 32'h140c8000, 32'h0, 32'hf0000000, 32'h1},{32'h0, 32'h0, 32'h0, 32'h316ad1c0, 32'h127a, 32'h0, 32'h2600000, 32'h0, 32'h980007c, 32'h3e02605c, 32'hb8, 32'h0, 32'ha0000000, 32'h0},{32'h0, 32'h0, 32'h0, 32'ha3385240, 32'h8d5, 32'h0, 32'h2e0c400, 32'hc40c000, 32'hc00002e, 32'h0, 32'h42000108, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h29ab41c0, 32'h1bbe, 32'h0, 32'h3000000, 32'h0, 32'h1e800000, 32'h420f4, 32'h42000000, 32'he0000, 32'hc8000380, 32'h0},{32'h0, 32'h0, 32'h0, 32'h27272340, 32'hc55, 32'h0, 32'h3a00000, 32'h1a800, 32'h1a832026, 32'h26000, 32'h7c0c81b0, 32'h1b0000, 32'hf00007c0, 32'h0},{32'h100, 32'h6000000, 32'h1c05000, 32'h5ee55a40, 32'hc61608d5, 32'he285e30f, 32'h710e543, 32'hd41c81b, 32'h1c81b072, 32'h2607406c, 32'h740001ac, 32'h881ac260, 32'h101c06b0, 32'h1},{32'h0, 32'h4014000, 32'h1c, 32'hd159c5a6, 32'hb71a49ca, 32'he2e5e50d, 32'h3007963, 32'hc813037, 32'h13040080, 32'h3806b000, 32'h730c81cc, 32'h641f8190, 32'hcc1f07e0, 32'h1},{32'h401c0, 32'h14000, 32'h18, 32'h76bd5de0, 32'hca96cdd2, 32'he3248a8a, 32'h4b09943, 32'hc1a43e, 32'h13033066, 32'h3e07d02c, 32'h4d088110, 32'hc8058340, 32'h90040680, 32'h1},{32'h180, 32'h401c000, 32'h0, 32'h62b441e5, 32'h6511a9be, 32'hce85dd49, 32'h7b0a8c3, 32'h1b800, 32'h1602d054, 32'h1c015088, 32'h44070194, 32'h158000, 32'h342b0380, 32'h1},{32'h70100, 32'h18000, 32'h5000, 32'hd5376ec0, 32'hca9b9153, 32'h3304e50f, 32'h6912093, 32'h15432, 32'h2402a000, 32'h7055028, 32'h7e01c150, 32'hfc1f4180, 32'h98000300, 32'h1},{32'h42800, 32'h70, 32'h0, 32'h60000006, 32'hea4f717d, 32'ha1446ace, 32'h86402d92, 32'hf40bc31, 32'h1f40b036, 32'h4d0360f4, 32'h321340c8, 32'h1c0580c0, 32'h5c070660, 32'h0},{32'h18000000, 32'h10070, 32'h0, 32'he7692d25, 32'had9db17d, 32'h4187ae88, 32'h8006ce3, 32'hc0d803, 32'h5440031, 32'h10065050, 32'h280401f8, 32'h54080000, 32'hf41507e0, 32'h1},{32'h14000000, 32'h18070, 32'h0, 32'h58f66f04, 32'hba9759bc, 32'hcd45824e, 32'h3a078e3, 32'h840c800, 32'h9c2107d, 32'h2f064, 32'h32068000, 32'h781901f0, 32'ha4320300, 32'h0},{32'h5010c, 32'h7000000, 32'h0, 32'h12bd0000, 32'h7c19eddb, 32'h71c59d4f, 32'h6305ea3, 32'h700c41c, 32'h1f821030, 32'h1038000, 32'h10c, 32'h10020010, 32'h1a0380, 32'h2},{32'h0, 32'h18050, 32'h4000, 32'h17250007, 32'hcb93316b, 32'ha136e54d, 32'h1400142, 32'h3c00000, 32'h1ec14082, 32'h4104303c, 32'h280781a0, 32'h2c0e41e0, 32'hcc010680, 32'h0},{32'h1c000000, 32'h50, 32'h18, 32'hf179af44, 32'h896c9c6, 32'hd5a47a8b, 32'h3c04ce3, 32'hd414000, 32'h19422027, 32'h28042074, 32'h7d0041a8, 32'h500e8010, 32'hf42303e0, 32'h0},{32'h40, 32'h3380060, 32'h1400008, 32'hf6ad0004, 32'h389f0f6a, 32'h2b24b0d, 32'h6b0e178, 32'hc817, 32'hdc39020, 32'h2684e040, 32'h6d09c1b4, 32'h68000000, 32'he4260450, 32'h0},{32'h1c000080, 32'hc000, 32'h4c4000, 32'h5, 32'h5939698, 32'hf1e99576, 32'h730dd8c, 32'h980f000, 32'hf017065, 32'h170750d4, 32'h4c08c1a8, 32'h660cc000, 32'hfc3806d0, 32'h0},{32'hc050000, 32'h7000000, 32'h1802000, 32'h28000004, 32'h179f958e, 32'h26ee06e6, 32'h4401db8, 32'h1c1f407, 32'h380f081, 32'hb04603c, 32'h46000114, 32'hac1fc000, 32'h240b0650, 32'h0},{32'h800004e, 32'h4018000, 32'h3014, 32'h679a5e80, 32'hc71a5ba5, 32'h8167e68d, 32'h4d0ab14, 32'hec15008, 32'h1d810067, 32'h45040, 32'h390e40e4, 32'h241a4070, 32'h58070560, 32'h1},{32'h8600000, 32'h4004050, 32'h0, 32'h52000000, 32'hcc91759b, 32'hdd58020b, 32'h640f947, 32'hb600000, 32'h15401059, 32'h3207105c, 32'h1000003c, 32'h4008000, 32'hc03e0100, 32'h0},{32'h14c000c0, 32'h4000000, 32'h1c00000, 32'h58000000, 32'h251dcbc5, 32'h81130ed2, 32'h910c5a8, 32'h6e19010, 32'hc81d07b, 32'h20004, 32'h3a04426c, 32'h44110010, 32'h100000f0, 32'h1},{32'h401c0, 32'h280010, 32'h3018, 32'h64c45000, 32'hf597936e, 32'h89c7aacc, 32'h3700d8d, 32'hc01c00, 32'h5c1e03c, 32'h108800cc, 32'h210f80cc, 32'h641e0, 32'hf8340000, 32'h1},{32'h0, 32'h0, 32'h8c4280, 32'haa000000, 32'h39953bbd, 32'h85a6e49e, 32'h420b887, 32'h640c01d, 32'h1f80407a, 32'h2e029010, 32'h3a0000c8, 32'h7a0fc328, 32'hd01c02b0, 32'h0},{32'h8000000, 32'h4018000, 32'h5000, 32'he0186840, 32'h989b759d, 32'h71181b93, 32'h14b, 32'hfc05800, 32'he01b043, 32'hb03901c, 32'h3101c00c, 32'h24000, 32'hf0190340, 32'h1},{32'h18020140, 32'h0, 32'h1c00000, 32'h4, 32'h389f1378, 32'h1490d2a, 32'h100174, 32'h13410c14, 32'hf84901f, 32'ha03c058, 32'h9a0280a0, 32'h58050000, 32'hc0a0170, 32'h0},{32'hc000000, 32'h82000000, 32'h14c0004, 32'hdcc4c820, 32'h3a97917d, 32'he686e2cb, 32'h6a00102, 32'h10020800, 32'ha43d083, 32'h1d08005c, 32'h3d0061a4, 32'h7e0e03e0, 32'hb02f0290, 32'h1},{32'h10001800, 32'h0, 32'h0, 32'h1, 32'h78b05a02, 32'hf315e49b, 32'h8720e099, 32'he41ac28, 32'h2104d021, 32'h390640f8, 32'h741341d0, 32'hd0000000, 32'h1c3a0740, 32'h1},{32'h22800, 32'h3004040, 32'h0, 32'h84910000, 32'ha76e157e, 32'hf172e5e2, 32'h83309949, 32'h381cc1e, 32'hbc0e010, 32'h804f020, 32'h80000d4, 32'h10040000, 32'h380900e0, 32'h1},{32'h1c013100, 32'h2180050, 32'h0, 32'hc2808000, 32'h3a9eee5e, 32'h25868b09, 32'h80f02d65, 32'h2c13407, 32'h7c0b00f, 32'h23814000, 32'h2407c1c4, 32'h0, 32'hc41e0180, 32'h1},{32'h0, 32'h1000640, 32'h805000, 32'hc0000000, 32'hc0001505, 32'hf3725389, 32'h8e0d0f4, 32'h841a021, 32'h8400002, 32'h3b01708e, 32'h5600015c, 32'h803c000, 32'he0000470, 32'h1},{32'h0, 32'h50, 32'hc81000, 32'h82208000, 32'hbd1399bb, 32'h723b458a, 32'h80011c, 32'h1c11024, 32'hc07077, 32'h24008000, 32'h300000c0, 32'h615c080, 32'h88080130, 32'h1},{32'h50000, 32'h10070, 32'h1308, 32'h6ae0c020, 32'hc89b3a92, 32'h8f06e20f, 32'h20000db, 32'h3c08404, 32'hcc2203e, 32'h3010, 32'h7f07c108, 32'h800c4228, 32'h9c2003c0, 32'h1},{32'h14000100, 32'h3000010, 32'h0, 32'h0, 32'hbd5c5998, 32'h71eab24a, 32'h706958, 32'hc800000, 32'hec3303d, 32'h3109a000, 32'h3c13408c, 32'h64000000, 32'h88000670, 32'h1},{32'h1400008e, 32'h18040, 32'h0, 32'h9e170000, 32'hc4162c4c, 32'hf2b71a0d, 32'h81087b5, 32'h4c04000, 32'h2400033, 32'h1d033070, 32'h120001fc, 32'h640a8000, 32'ha8000340, 32'h0},{32'hc0, 32'h10000, 32'h0, 32'h0, 32'h2c11cf48, 32'hb14b0c66, 32'h5d11c8b, 32'h1201f835, 32'h1f01f032, 32'hf02c, 32'h4a000128, 32'hcc2041f0, 32'h83306c0, 32'h0},{32'h14020000, 32'h401c000, 32'h1300, 32'hd2ac8e60, 32'hcda2f072, 32'h36e55b, 32'h6c0018a, 32'h100e436, 32'h9b, 32'h403d010, 32'h6c000054, 32'hd40a8, 32'hb8380080, 32'h1},{32'h900, 32'h8000, 32'h28000000, 32'he6000003, 32'h84939155, 32'h69c5e64a, 32'h86b0e992, 32'h6c0a41f, 32'he80003a, 32'h1c02d000, 32'h820000e8, 32'h81901d0, 32'h54368761, 32'h2},{32'h800004a, 32'hc040, 32'h0, 32'h6, 32'hb846c000, 32'hd3665398, 32'h830e6db, 32'hcc1f031, 32'h26c42081, 32'h2b03b128, 32'h198, 32'hc2502b0, 32'hd42605f1, 32'h1},{32'h140, 32'h83000000, 32'h800004, 32'h6, 32'h30001168, 32'h2e19bb13, 32'h4d0015c, 32'h300600e, 32'h6000085, 32'h701c000, 32'h690121d4, 32'h20038130, 32'h3c130750, 32'h1},{32'hca00000, 32'h8040, 32'h0, 32'h0, 32'h19472d48, 32'h5e85c2d8, 32'h6a0e542, 32'h2e1c800, 32'h5c2b01d, 32'h3a0110e8, 32'h480d81b0, 32'h0, 32'h4c2c0740, 32'h0},{32'h40000, 32'h118000, 32'h400014, 32'h0, 32'h97138ac0, 32'hcdfa854c, 32'h11d, 32'h10c1a, 32'h4000000, 32'h12857000, 32'h570000fc, 32'hbc0d8080, 32'h190, 32'h0},{32'hc000100, 32'h7000000, 32'h28800018, 32'h1, 32'hc6968000, 32'h732762cf, 32'h9084b3, 32'h3c07800, 32'h5819099, 32'h1a077020, 32'h310900c4, 32'h300601a0, 32'he4088050, 32'h1},{32'h40000, 32'h0, 32'h1100, 32'h0, 32'hc7ec7300, 32'hf1b58ae8, 32'h18b, 32'h244d, 32'h28000000, 32'h40000, 32'h110000f8, 32'h2811c318, 32'h700a0a00, 32'h2},{32'h0, 32'h6014000, 32'h80400c, 32'h6338ad20, 32'h8512968d, 32'h646e64a, 32'h103, 32'h11c0d050, 32'h23800045, 32'h4709b11c, 32'h230600f4, 32'h400044d0, 32'hc0360411, 32'h1},{32'h0, 32'h3000000, 32'h800010, 32'he2000001, 32'h9b91b48c, 32'hf30f02c9, 32'h6200084, 32'h1b033, 32'h6c, 32'h33018000, 32'h10d818c, 32'h301b8000, 32'ha4000630, 32'h1},{32'h23800, 32'h64000000, 32'h14c0004, 32'h0, 32'h959e4000, 32'h5b066475, 32'h888070f3, 32'hec0b, 32'he000036, 32'h1f03c000, 32'h3502612c, 32'hda0ac050, 32'h28460670, 32'h0},{32'hca00000, 32'h4000010, 32'h0, 32'h0, 32'hdd112000, 32'h6e32120a, 32'h7c0f54b, 32'h121f000, 32'hd43a091, 32'h3a07e000, 32'h68000024, 32'hfc1f8340, 32'h43a0660, 32'h2},{32'h0, 32'h4000, 32'hc00000, 32'h2, 32'hc8a6a000, 32'h49aa76b6, 32'h6d0acbc, 32'hb400000, 32'h15800064, 32'h4106d000, 32'h380000e8, 32'h0, 32'hbc2e0710, 32'h1},{32'hc000000, 32'h4000000, 32'h400000, 32'h0, 32'h2b912000, 32'h6e0e046c, 32'h660e542, 32'hec1d800, 32'h1983203b, 32'h38000000, 32'h15c, 32'hd8000000, 32'hc0000770, 32'h1},{32'h4000000, 32'h8000, 32'h4000, 32'h0, 32'h80000000, 32'he90b8df7, 32'h740014a, 32'he805807, 32'h600e067, 32'h95000, 32'h100001d0, 32'h9c3b0, 32'h68000870, 32'h0},{32'h10000, 32'h0, 32'h1000000, 32'h9c000000, 32'h8ae46b48, 32'h5f446d30, 32'h740e502, 32'hac0643a, 32'h1b02b019, 32'h1406c050, 32'h56000120, 32'h88000000, 32'hd8140750, 32'h1},{32'h0, 32'h1000000, 32'h0, 32'h3900002, 32'h882c720d, 32'hceaebeb6, 32'h3401d14, 32'h8810840, 32'h2003e012, 32'h9075000, 32'h100001b4, 32'hc8000, 32'h64230000, 32'h1},{32'h0, 32'h10000, 32'h8, 32'h0, 32'h18eec370, 32'he6f84e98, 32'h320014a, 32'h0, 32'h6800000, 32'h18011000, 32'h5f00c060, 32'h17c0e0, 32'h78030000, 32'h0},{32'h10030000, 32'h18050, 32'h1c02000, 32'h0, 32'hc499f010, 32'h86876a0f, 32'h4a001a8, 32'h781244c, 32'h420001, 32'h107c, 32'h4e000138, 32'h64000, 32'h841f0150, 32'h0},{32'h0, 32'h14032, 32'h0, 32'h2, 32'h1c978000, 32'h42770552, 32'h76000ed, 32'hec1f83e, 32'h2844789a, 32'h2808f0a0, 32'h4c100280, 32'h0, 32'h743a0000, 32'h2},{32'h0, 32'h0, 32'h400180, 32'h0, 32'ha8584000, 32'hbe2e9dd3, 32'h7e0f58c, 32'hb000000, 32'h1d80007e, 32'h39066000, 32'h560001b0, 32'hc81c44d8, 32'he0000370, 32'h1},{32'h0, 32'hc000, 32'h1000, 32'h0, 32'ha92c4080, 32'h729145b7, 32'h80c977, 32'h9800000, 32'h19000038, 32'h19000, 32'h38000130, 32'h4c1bc330, 32'h281304e0, 32'h2},{32'h40, 32'h0, 32'h2000, 32'h0, 32'h4686b48, 32'h36f0559c, 32'h3f065ba, 32'hf81f800, 32'h64, 32'h740d0, 32'h34060000, 32'h2c3e0, 32'hf8000681, 32'h1},{32'h0, 32'h0, 32'h4, 32'h0, 32'h255a6390, 32'haf6f721a, 32'h4e0998b, 32'h2c20800, 32'h7a, 32'h3207f104, 32'h69030208, 32'h0, 32'h40000180, 32'h1},{32'h0, 32'h10, 32'h0, 32'h3, 32'h8c584000, 32'hcd577eb6, 32'h570c908, 32'h3800, 32'hec00064, 32'h4e018000, 32'h9c0cc048, 32'h2800c0, 32'h74000a00, 32'h1},{32'h20000, 32'h1280000, 32'h1000000, 32'h0, 32'hc7123268, 32'h3e18e288, 32'h670d9bb, 32'h1dc0d, 32'h1e00001a, 32'h886e0e8, 32'h6e0f01c4, 32'hdc000000, 32'h58000010, 32'h0},{32'h33000, 32'h10050, 32'h1000, 32'h2, 32'h279a8098, 32'h67655b8b, 32'h85600164, 32'hb40743a, 32'h1b414028, 32'h6d0b8, 32'h56070170, 32'h1dc1c0, 32'h6c2c0000, 32'h0},{32'h4000000, 32'h640, 32'h0, 32'h83602422, 32'hc0001506, 32'hf20d9ddd, 32'h1800107, 32'h3011000, 32'h4417057, 32'h29092, 32'h1a000000, 32'h34000000, 32'hdc180440, 32'h1},{32'hc000000, 32'h4000000, 32'h2000, 32'h0, 32'ha591c000, 32'hf30a0dc9, 32'h9a, 32'h342043a, 32'h13, 32'h101c01c, 32'h76000064, 32'hc0dc0f0, 32'hd8000160, 32'h1},{32'h0, 32'h0, 32'h800000, 32'h0, 32'hd5c46000, 32'hbaea0ca6, 32'h4009c8c, 32'h15800, 32'h1381f056, 32'h40078, 32'hd4, 32'ha0000000, 32'h381f01f0, 32'h1},{32'h8000000, 32'h0, 32'hc00000, 32'h0, 32'h194f58b0, 32'h2c08a552, 32'h4c0d9b4, 32'ha00a000, 32'h1b828041, 32'h6c050, 32'h6e00013c, 32'h0, 32'h383709b0, 32'h1},{32'h10030080, 32'h4000, 32'h0, 32'h0, 32'h50a2f898, 32'h25c4a075, 32'h770a9b9, 32'hec2843f, 32'h1603606d, 32'h510f8, 32'h810e0000, 32'he0000000, 32'h68000740, 32'h1},{32'h1800, 32'h0, 32'h1000000, 32'h0, 32'h1a6d0000, 32'hbf3315d4, 32'h86c000ba, 32'h16433, 32'h6c, 32'h3706c000, 32'h780dc1e0, 32'he01c0370, 32'h98000270, 32'h1},{32'h80, 32'h40, 32'h400000, 32'h3, 32'h17120040, 32'h357263e5, 32'h39021ab, 32'h1c00000, 32'h1d41006c, 32'h320fc, 32'h7e0441c0, 32'he00d0110, 32'h340904f0, 32'h2},{32'h0, 32'hc000, 32'h2000, 32'hc4000000, 32'h6482e14, 32'hbf774aed, 32'h76098da, 32'h1d800, 32'h2083a000, 32'h6909c, 32'h82000138, 32'hc81fc000, 32'h810, 32'h0},{32'h0, 32'h800, 32'hc00004, 32'h2, 32'ha0000000, 32'hd21b9e2b, 32'h38084e5, 32'h441301c, 32'h8800044, 32'h83032, 32'h190401f8, 32'h9c1f8230, 32'h44330850, 32'h1},{32'h10000000, 32'h3000010, 32'h2000, 32'h18bc0120, 32'h1acc, 32'hdedb6800, 32'h147, 32'h5400000, 32'h4c15075, 32'h2c000000, 32'h58054274, 32'h54284000, 32'h580, 32'h0},{32'h18000140, 32'h8032, 32'h400000, 32'h7, 32'h751e2000, 32'hb9667d49, 32'h57000a2, 32'he806c2e, 32'h1e414829, 32'h1c06f0f0, 32'h78000170, 32'h1d8000, 32'h643b06f0, 32'h1},{32'h20000, 32'h4000, 32'h0, 32'h0, 32'hc0000000, 32'he5d79a6e, 32'h4400108, 32'h16c00, 32'h1743a038, 32'h1c05d070, 32'h18000110, 32'h740c00c0, 32'hd81d0760, 32'h1},{32'h80, 32'h0, 32'hc, 32'h18000000, 32'had402e68, 32'haed14a2a, 32'h190b169, 32'h16033, 32'h7033000, 32'h64000, 32'h1b000000, 32'h160000, 32'h40000580, 32'h0},{32'h40000, 32'h60000000, 32'h1000, 32'h0, 32'hba204000, 32'h65446609, 32'h3e05559, 32'h15c00, 32'ha82000e, 32'h9012000, 32'h7700e0a8, 32'h741f0, 32'h2a0, 32'h0},{32'h8040000, 32'h10, 32'h0, 32'h0, 32'hbab47a10, 32'h49448509, 32'h340951b, 32'h2c0a40d, 32'h13c0b03f, 32'h0, 32'h250, 32'hdc250000, 32'hd8190510, 32'h0},{32'hc000000, 32'h11, 32'h0, 32'h0, 32'hcd250b00, 32'hc337e66b, 32'h1001ccd, 32'he81d83a, 32'h1bc28851, 32'h0, 32'h0, 32'h580b0090, 32'hbc140780, 32'h1},{32'h40, 32'h0, 32'h4000, 32'h3, 32'hac5c4000, 32'hb5696632, 32'h7f109ad, 32'h2101e, 32'h2103e07c, 32'h0, 32'h71000000, 32'h19c200, 32'h6c200000, 32'h1},{32'h0, 32'h2194000, 32'h90, 32'h0, 32'h80000000, 32'h6d396d2b, 32'h200214b, 32'h11c0f81e, 32'hd00f090, 32'h3c87f07c, 32'h7f0241bc, 32'h1bc388, 32'h40000000, 32'h0},{32'h0, 32'h62000000, 32'h0, 32'h1, 32'hc9e71418, 32'h5b687eab, 32'h4e03d75, 32'hb01380f, 32'h1380f04e, 32'h27056000, 32'h2306a1c4, 32'h140370, 32'h4c370000, 32'h0},{32'h88, 32'h5004000, 32'h180001c, 32'h3808000, 32'h6d198d4d, 32'h7335dc4d, 32'h7707379, 32'h10408840, 32'h20c11080, 32'h1004f104, 32'h670fc1fc, 32'h198000, 32'h4f0, 32'h0},{32'h0, 32'h0, 32'h1000, 32'h0, 32'h80000000, 32'h5ecfcd63, 32'h7e00136, 32'h500a800, 32'ha814023, 32'h1a000000, 32'h7e0681f8, 32'h5411c150, 32'h800, 32'h2},{32'h8000000, 32'h23000000, 32'h0, 32'h0, 32'h8a5f1178, 32'hb750569c, 32'h320bcba, 32'hd000, 32'hb80002b, 32'h0, 32'h59056164, 32'h68000, 32'h780001a0, 32'h1},{32'h0, 32'h4a00, 32'h2010, 32'h0, 32'hc4536000, 32'h3345e60b, 32'h80000a2, 32'hb01741c, 32'h2000080, 32'h2b079062, 32'h190ec1f8, 32'h141dc230, 32'h68050460, 32'h1},{32'h0, 32'h0, 32'h800000, 32'h86d18723, 32'ha0000f12, 32'h2ef145a1, 32'h660009a, 32'hcc00000, 32'h404101c, 32'h410580c8, 32'h580cc160, 32'h76198000, 32'h1c340770, 32'h1},{32'h88, 32'h0, 32'h1000, 32'h3208000, 32'hab506e0c, 32'ha633add9, 32'h5907f77, 32'h19c09, 32'h18, 32'h18104, 32'h66000048, 32'h81643b0, 32'h400d0761, 32'h0},{32'h86, 32'h1000000, 32'h1000000, 32'h0, 32'h90000d50, 32'h666e5da4, 32'h2b08304, 32'h3006000, 32'h32, 32'hc013000, 32'h180000ac, 32'h38000000, 32'h6f0, 32'h0},{32'h80, 32'h0, 32'h0, 32'h3, 32'hc1456000, 32'h604e08ed, 32'h1b00177, 32'he000, 32'ha000028, 32'h16010000, 32'h2c0e0254, 32'h741c0000, 32'hdc0906e0, 32'h0},{32'h0, 32'h0, 32'h801000, 32'h3, 32'h14c80bc0, 32'h3c34706d, 32'hc5, 32'h0, 32'h84, 32'h3706e000, 32'h7e0001f8, 32'hdc0b42f0, 32'he4000790, 32'h1},{32'h0, 32'h40, 32'h1000, 32'h0, 32'h6938000, 32'hcace15a0, 32'h5000115, 32'h0, 32'hd42803e, 32'h52000, 32'h500a4000, 32'h104290, 32'h40000000, 32'h1},{32'h60000, 32'h50, 32'h4004, 32'h2, 32'ha69a43b0, 32'h39a57d4d, 32'h7e0e083, 32'hcc13c33, 32'h13c4b091, 32'h4e0fc, 32'h13100258, 32'hcc1bc000, 32'h8c100200, 32'h0},{32'h40, 32'h0, 32'h3000, 32'h42a08000, 32'h90000292, 32'hd7537dd7, 32'h1f0ad0d, 32'h1f02d, 32'h20037000, 32'h0, 32'h1b8, 32'h4144370, 32'h700005b1, 32'h1},{32'h11000, 32'h4000000, 32'h0, 32'h0, 32'h50000000, 32'ha2985c1b, 32'h8880019d, 32'ha020411, 32'h13828083, 32'h1502a064, 32'h2a0100d4, 32'h6c200000, 32'h401b0500, 32'h1},{32'h30000, 32'h0, 32'h0, 32'h4e04402, 32'hb4514113, 32'hf2b4ba66, 32'h1a7, 32'hac00, 32'h12019046, 32'hd048030, 32'h34000118, 32'hac1b0, 32'h41b01a0, 32'h2},{32'hc0, 32'h80000000, 32'h1400308, 32'h7, 32'h654e2170, 32'hb645a40d, 32'h5f0ac9a, 32'h16000, 32'h1682a000, 32'h60000, 32'h370ee000, 32'hb806c238, 32'hec000470, 32'h0},{32'h80, 32'h5018000, 32'h10, 32'h0, 32'hb9178000, 32'h8644e52a, 32'h810b58d, 32'h1682b, 32'h1e000000, 32'h3c059104, 32'h590ec164, 32'hcc050000, 32'h780000b0, 32'h0},{32'h80, 32'h0, 32'h4000, 32'h0, 32'h14306000, 32'hee2fa4d6, 32'h670ed8c, 32'h0, 32'h4000000, 32'h1a01208c, 32'h760bc118, 32'h8c1dc2f0, 32'ha4000780, 32'h1},{32'h0, 32'h0, 32'h400000, 32'h2, 32'ha9500000, 32'hbe0b9edc, 32'h18070d8, 32'h14000, 32'he80003a, 32'h50074, 32'h1c0, 32'h9c1c0370, 32'h6c1d0850, 32'h0},{32'h0, 32'h2000000, 32'hc80000, 32'h1, 32'h86361a00, 32'hda7ba497, 32'h7600134, 32'h6405, 32'h1780400a, 32'h3c0780bc, 32'hdc, 32'h761d81c0, 32'h743c01d0, 32'h0},{32'h0, 32'h22000000, 32'h3000, 32'h0, 32'h2d312000, 32'he66da459, 32'h380016a, 32'h201000c, 32'h1002e06e, 32'h5c000, 32'h7105a0b4, 32'h2404c070, 32'h680003e0, 32'h0},{32'h12080, 32'h0, 32'h0, 32'h80000003, 32'hb00008cd, 32'h568ac5da, 32'h8850012d, 32'h2141f, 32'h9000000, 32'h2606f000, 32'h94000148, 32'h148120, 32'h84110000, 32'h1},{32'h10000080, 32'h2000c000, 32'h1800000, 32'h5, 32'h47478000, 32'h4126e34d, 32'h510ccc2, 32'h380e80e, 32'h4f, 32'h8053074, 32'h510a61a0, 32'h741a0330, 32'h84340210, 32'h0},{32'h20000, 32'h0, 32'h4, 32'h44000000, 32'h1b12, 32'he66bc31b, 32'h8205978, 32'h19c40, 32'h25c00080, 32'h6e0fc, 32'h81000000, 32'h14028000, 32'h2e0, 32'h0},{32'h0, 32'h7000000, 32'h1005018, 32'ha4000000, 32'h1d9d4c58, 32'hf344e5a6, 32'h360b192, 32'hbc00000, 32'h4e, 32'h2f058000, 32'h2b0a00ac, 32'hc4204280, 32'h74280810, 32'h1},{32'h4000000, 32'h10000, 32'h860000, 32'h0, 32'hd5938f18, 32'h723aba6c, 32'h2a121b9, 32'h5421048, 32'h51, 32'h150350d0, 32'h800cc22c, 32'ha21a0400, 32'hb0370, 32'h2},{32'h8000000, 32'h3000010, 32'h0, 32'h0, 32'ha63e6e40, 32'hef0de5e3, 32'h5810194, 32'hb42001f, 32'h12400047, 32'h56000, 32'h5800006c, 32'h800dc200, 32'h800, 32'h0},{32'hc000000, 32'h10, 32'h0, 32'h0, 32'hbc84000, 32'hb70ade9c, 32'h82000bc, 32'h540a800, 32'h18400061, 32'h58000, 32'h2a0000d0, 32'h80d8400, 32'h361, 32'h0},{32'h0, 32'h11, 32'h3000, 32'h0, 32'hc04b8000, 32'haeeec2a0, 32'h5b109a6, 32'h21000, 32'h1e441846, 32'h34054, 32'h2206c000, 32'h6c07c150, 32'h88100800, 32'h0},{32'h30100, 32'h4000, 32'h800000, 32'h82000000, 32'he000136d, 32'h3f0ada12, 32'h1907cb9, 32'h4004c00, 32'h1400904e, 32'h8047024, 32'h5f080088, 32'h80088000, 32'h790, 32'h0},{32'h0, 32'h3000010, 32'h0, 32'h0, 32'hfa584008, 32'hd59782f6, 32'h600138, 32'h1e02f, 32'hec00000, 32'h1c05e014, 32'h700001c4, 32'h1e8000, 32'h30000000, 32'h0},{32'h14000000, 32'h8010, 32'h20000000, 32'h3, 32'h99e90000, 32'hf30564a3, 32'h10030e2, 32'h2c07, 32'h17c2306f, 32'h407908c, 32'h1a1200d0, 32'h68310, 32'he40d8620, 32'h1},{32'h10000, 32'h0, 32'h0, 32'h0, 32'hed645598, 32'hf1506b36, 32'h5a000f8, 32'h10410, 32'h1741a000, 32'h0, 32'h240b00d8, 32'h88000, 32'h70000360, 32'h1},{32'hc000100, 32'h0, 32'h0, 32'h5, 32'h17644000, 32'hc34f4332, 32'h67014aa, 32'h1e003, 32'he806095, 32'hd00a000, 32'hc00014c, 32'h68000, 32'ha40d0000, 32'h1},{32'h0, 32'h2000050, 32'h4000, 32'h0, 32'hb766a1a0, 32'hc705e4b3, 32'h66030c4, 32'h742c, 32'h1bc41082, 32'h16000000, 32'h2c0541a4, 32'h3802c000, 32'h600e05a0, 32'h1},{32'h0, 32'h0, 32'h8860010, 32'h0, 32'haaeac000, 32'hadcf8e50, 32'h820009d, 32'h1001f, 32'h6800040, 32'h5e000, 32'h51070000, 32'h5e050000, 32'hc428830, 32'h2},{32'h0, 32'h80000000, 32'h10c, 32'h0, 32'h1d138000, 32'h72d9c49e, 32'h4007d46, 32'h8024000, 32'h2400a016, 32'h0, 32'h63102000, 32'h16c288, 32'h48000160, 32'h2},{32'h4, 32'hc000, 32'h0, 32'h1, 32'hcc2b8000, 32'hea95402d, 32'h910577d, 32'h16800, 32'h1b800084, 32'h380690fc, 32'h5a0e0100, 32'hc168280, 32'h1c2c0501, 32'h2},{32'h40, 32'h0, 32'h0, 32'hc13842, 32'h30000d54, 32'hadf48e12, 32'h8105569, 32'h11800, 32'h20816000, 32'h68000, 32'h2c0d0000, 32'h104000, 32'h6c340000, 32'h1},{32'h14010000, 32'h10000, 32'h2180, 32'h0, 32'hc712bb08, 32'hca89060b, 32'h660b8f4, 32'h12c0ac40, 32'h47, 32'h4b02b0b8, 32'h681001a0, 32'h740dc2e8, 32'hc8000820, 32'h1},{32'h10000040, 32'h40000000, 32'h0, 32'h0, 32'ha76a0000, 32'h5e6bde5e, 32'h8501114, 32'ha02e, 32'hd00003b, 32'h502c0b8, 32'h37046188, 32'h100160, 32'he8050620, 32'h0},{32'h30000, 32'h1000000, 32'h0, 32'h0, 32'h96e24260, 32'hc55484d1, 32'h460a09d, 32'h2414423, 32'h4c24050, 32'h12020, 32'h5006c08c, 32'hd8000, 32'h0, 32'h0},{32'h20000, 32'h2, 32'h1000, 32'h3, 32'haa938f60, 32'hdecede49, 32'h600129, 32'h17c24, 32'h1c42380c, 32'h1101a090, 32'h22018040, 32'h1ec230, 32'h34090000, 32'h0},{32'h0, 32'h0, 32'h1008, 32'h84000000, 32'h30001174, 32'h5a6dca60, 32'h5e004fd, 32'h417800, 32'h2642f02a, 32'h30054, 32'h1b044008, 32'h18c1b0, 32'he81605e0, 32'h0},{32'h40000, 32'h30, 32'h0, 32'h9e000001, 32'haaa30068, 32'h6ed34aa5, 32'h2c00178, 32'hec00, 32'h9405008, 32'h39096000, 32'h1a054030, 32'h20000, 32'h74170000, 32'h1},{32'h40, 32'h0, 32'h0, 32'h0, 32'h28586070, 32'hf34f4d58, 32'h790b128, 32'h680b, 32'h25800000, 32'h12096000, 32'h72000160, 32'h70120, 32'h80000000, 32'h0},{32'hc000000, 32'h1000000, 32'h0, 32'h0, 32'h4dc04000, 32'h4719649d, 32'h38000d4, 32'h0, 32'h17804083, 32'h6052018, 32'h520a00b4, 32'h14000000, 32'h280001d1, 32'h2},{32'h10000, 32'h0, 32'h3000, 32'h0, 32'h2a684000, 32'hae359b9f, 32'h900008a, 32'h10430, 32'h5800052, 32'h600b0, 32'h1d000000, 32'h2142a0, 32'h70000000, 32'h1},{32'h0, 32'he5000000, 32'h80430c, 32'h0, 32'h194f2000, 32'hb507e6a8, 32'h410b562, 32'h4c24800, 32'h1c013092, 32'h2c070124, 32'h930b6104, 32'h1442d8, 32'h930, 32'h0},{32'h100, 32'h1000000, 32'h0, 32'h2000000, 32'h2000120d, 32'he275b6e2, 32'h2b0593b, 32'h14000, 32'h4000050, 32'h2902a000, 32'h520241c4, 32'h140170, 32'h48000870, 32'h0},{32'h0, 32'h30, 32'h400000, 32'h2, 32'h1b330000, 32'h35147b99, 32'h1b9, 32'h4010042, 32'hb434052, 32'h69048, 32'h80048100, 32'hc000000, 32'h24000851, 32'h1},{32'h40, 32'h3000000, 32'h800010, 32'h0, 32'hcb139518, 32'hcf2e5e21, 32'h5d10cfb, 32'h7400000, 32'h17000097, 32'h15000000, 32'h410581a4, 32'h141702d0, 32'h70000830, 32'h1},{32'h0, 32'h1000000, 32'h10, 32'h0, 32'h3a5c4058, 32'hf10d63e2, 32'h400b9b6, 32'h1001d, 32'h2182e000, 32'h340880d0, 32'h3708018c, 32'h38000000, 32'h20000480, 32'h1},{32'h600044, 32'h4014000, 32'h0, 32'h4a10000, 32'hca16538a, 32'hef0fd2cb, 32'h5108f5c, 32'h920204d, 32'h26800013, 32'h601b014, 32'h6206c08c, 32'h18048310, 32'h200009c0, 32'h0},{32'h10000, 32'h4014000, 32'h800000, 32'h0, 32'he8e00c10, 32'h2f34535e, 32'h1c01d34, 32'h12415, 32'h2180e000, 32'h4a023068, 32'h940980dc, 32'h178000, 32'h130, 32'h0},{32'h30000, 32'h4000000, 32'h0, 32'h0, 32'h2a1381c8, 32'he9cf8b26, 32'h31115d, 32'h1017c04, 32'ha, 32'h1b000000, 32'h5e01406c, 32'h228040, 32'h80050000, 32'h1},{32'h0, 32'h30, 32'h0, 32'h1, 32'h8b5c4000, 32'hb1397ba2, 32'h97035b6, 32'h8c08824, 32'h3424022, 32'h2018008, 32'h2000088, 32'h0, 32'hbc2d0000, 32'h0},{32'h0, 32'h20, 32'h0, 32'h0, 32'h8dc82348, 32'h4eb7cda1, 32'hc01117, 32'h1402001, 32'h25c00002, 32'h6000000, 32'h8a004094, 32'h0, 32'h28060000, 32'h2},{32'hc000000, 32'h4400, 32'h0, 32'h0, 32'ha461c000, 32'h26cfcc77, 32'h780e57c, 32'h12c00000, 32'h1804b05f, 32'hd0a6, 32'h60, 32'h168000, 32'h8b0, 32'h0},{32'h0, 32'h10050, 32'h4, 32'h2, 32'h31438000, 32'hdf44e518, 32'h900015d, 32'h741780b, 32'h1c44905e, 32'h1b071000, 32'h5d124188, 32'h154310, 32'h4c140000, 32'h2},{32'h0, 32'h0, 32'h800000, 32'h0, 32'h8aa42000, 32'hbdb185af, 32'h500f1ac, 32'h24c00, 32'h1c000082, 32'h760e0, 32'h0, 32'h241e8000, 32'h483c05d0, 32'h1},{32'h30000, 32'h2000040, 32'h0, 32'h6158000, 32'h9b139a1a, 32'h3254e4a6, 32'h2a045ba, 32'h14400, 32'h1a405022, 32'h4022000, 32'h14c, 32'hbc060, 32'hb80002e0, 32'h0},{32'h30000, 32'h4000000, 32'h440000, 32'h0, 32'ha0000000, 32'hb6d2da34, 32'h2a00158, 32'h14c00, 32'h25800048, 32'h16025000, 32'h2c, 32'h86220000, 32'hd0000870, 32'h1},{32'h30000, 32'h10000, 32'hc1000, 32'h5, 32'hc6138000, 32'h723a158d, 32'h8600144, 32'h17400, 32'h18000004, 32'h11069048, 32'h5a000090, 32'h92174020, 32'h24210890, 32'h1},{32'h2, 32'h2000000, 32'h4000, 32'h0, 32'h3d386908, 32'hda8ee423, 32'h5d082da, 32'h0, 32'h2806082, 32'h2d068018, 32'h8000074, 32'h4c050, 32'h20000840, 32'h1},{32'hc000000, 32'h0, 32'h400008, 32'h4, 32'haa380000, 32'hd628e5a4, 32'h9600136, 32'h3800000, 32'h2581200d, 32'h10044, 32'h63000090, 32'he8000000, 32'hb42709d0, 32'h0},{32'hc000080, 32'h1000000, 32'h0, 32'h0, 32'ha78000, 32'hd68bd5e4, 32'h5f10d09, 32'h1002800, 32'hb000087, 32'h16000000, 32'h254, 32'h28000, 32'h281600a0, 32'h2},{32'h0, 32'h0, 32'h1000000, 32'h2, 32'h345c0150, 32'hd364e618, 32'h400114, 32'h2400000, 32'h1009048, 32'h0, 32'h4000000, 32'h4010090, 32'h842405b0, 32'h1},{32'h20000, 32'h0, 32'h3000, 32'h0, 32'h472f4000, 32'hdec90b25, 32'h208156, 32'h8c50, 32'h2784709e, 32'h4d005018, 32'ha0000028, 32'h84074170, 32'hb8160040, 32'h0},{32'h10000, 32'h0, 32'hc, 32'h82a08000, 32'hd9c04bde, 32'he691b212, 32'h4c000ea, 32'hc3a, 32'h2, 32'h4a094004, 32'h8b000168, 32'h90000000, 32'h340205c0, 32'h0},{32'h20000, 32'h0, 32'h3000, 32'h1, 32'ha0678000, 32'ha63a9416, 32'h5e00169, 32'h5018400, 32'h97, 32'h0, 32'h5e06c148, 32'h24c000, 32'hec2a0000, 32'h1},{32'hc020100, 32'hc1000000, 32'h0, 32'h5, 32'hc1df8000, 32'hea05e249, 32'h5100ce7, 32'hc017c11, 32'h1804e093, 32'h4d09c120, 32'h9302618c, 32'hb4240000, 32'h4c120780, 32'h1},{32'h0, 32'h0, 32'hc, 32'h84110002, 32'h700009ca, 32'hce51ad17, 32'h80a0cd, 32'h12808809, 32'h480000a, 32'h4a052000, 32'h85024148, 32'h1ec000, 32'he40004e0, 32'h1},{32'h0, 32'h0, 32'h800000, 32'h0, 32'h2b6801c0, 32'h5e8fcc37, 32'h115, 32'h12c1480e, 32'h1d00002c, 32'h0, 32'h12000000, 32'h94078000, 32'h280002f0, 32'h1},{32'h80, 32'h4000, 32'hc, 32'h4, 32'hc4117608, 32'h32f40609, 32'h4900197, 32'h24800, 32'h1a014092, 32'h2d004, 32'h89030010, 32'h220000, 32'hc490920, 32'h1},{32'h40, 32'h8000, 32'h0, 32'h0, 32'h384c0000, 32'haad5c328, 32'h6113497, 32'h304d, 32'h0, 32'h46025118, 32'hc004268, 32'h18000, 32'h20000060, 32'h0},{32'h0, 32'h4000, 32'h860000, 32'h0, 32'hc7230000, 32'hcf30da9e, 32'h117, 32'he807000, 32'h3446096, 32'h5b000, 32'h8c000000, 32'h1a0482a0, 32'h50290850, 32'h1},{32'h80000000, 32'h1, 32'h10, 32'h0, 32'h2b5c2000, 32'h55096e18, 32'hed, 32'h0, 32'h944a88c, 32'h2c004, 32'hb000230, 32'h180280e0, 32'h700d08a0, 32'h0},{32'h80, 32'h0, 32'h0, 32'hc4000001, 32'h30000092, 32'hd9096a98, 32'hb09109, 32'h0, 32'h80300c, 32'hc000, 32'ha000010, 32'h0, 32'h24250060, 32'h2},{32'h10140, 32'h20, 32'h10c0000, 32'h0, 32'h54939b08, 32'h5a141aa9, 32'h300127, 32'h1381244f, 32'h144f013, 32'h9a030, 32'h92138000, 32'ha000000, 32'h48000430, 32'h2},{32'h40000c0, 32'h0, 32'h2000, 32'h0, 32'he0000000, 32'h65ecba26, 32'hd02559, 32'h2428401, 32'h2800009f, 32'h5009a000, 32'h8a014028, 32'h140bc000, 32'h704605a1, 32'h1},{32'h0, 32'h4000, 32'h0, 32'h32000003, 32'he4285bb8, 32'h51704ade, 32'h119, 32'h1800, 32'h1000078, 32'h950f0, 32'h4000240, 32'h240000, 32'h643d07a0, 32'h2},{32'h6, 32'h10, 32'h8a6000, 32'h4, 32'h64954000, 32'h41daa4cd, 32'h5f126cc, 32'h27005, 32'h14c4d000, 32'h4d09c140, 32'ha000280, 32'hf21e4000, 32'h94060550, 32'h0},{32'h8000100, 32'h10, 32'h0, 32'h0, 32'h90000000, 32'he2119e5c, 32'h230bd2a, 32'h2402800, 32'h27429061, 32'h2f091000, 32'h28, 32'h1e83c0, 32'he81c02e0, 32'h1},{32'h800000, 32'h8000, 32'h0, 32'h6e000000, 32'hcc407510, 32'hed0d6289, 32'h2200114, 32'h5a18000, 32'h1e000095, 32'h530f0, 32'h18, 32'hc0000000, 32'h90030780, 32'h0},{32'h10080, 32'h0, 32'hc00000, 32'h0, 32'hc9aa8000, 32'hc168c2f5, 32'h530449a, 32'h25c14, 32'h9000092, 32'h2a048, 32'h0, 32'h7c000, 32'h904a04b0, 32'h0},{32'hc010000, 32'h8000, 32'h0, 32'h0, 32'h40cb8000, 32'ha668e4f7, 32'h16c, 32'h24c4b, 32'h25027005, 32'h89128, 32'h7602c050, 32'h38058000, 32'h704c0931, 32'h2},{32'h30040, 32'h0, 32'h2000, 32'hc2000000, 32'h9000080a, 32'h3e75a65c, 32'h9b000c8, 32'h9c03429, 32'h94, 32'h108d128, 32'h60000230, 32'h1c000, 32'h420, 32'h0},{32'h86, 32'h40, 32'h1400000, 32'h0, 32'hc8440000, 32'hdb2a0b89, 32'h1d12f3b, 32'h13847, 32'hb400000, 32'h94000, 32'h68, 32'h38128000, 32'h400000d0, 32'h2},{32'h100, 32'h0, 32'h2000, 32'h0, 32'h16138000, 32'ha258e2e0, 32'h4912599, 32'h24847, 32'h8d, 32'h4000, 32'h4a054000, 32'h2022c030, 32'h41, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h16a84370, 32'h2f0fdc94, 32'h1c12d9a, 32'h25800, 32'hd, 32'h9c134, 32'h0, 32'h1d8000, 32'h68000920, 32'h0},{32'h100, 32'h0, 32'h0, 32'h5, 32'h294c2000, 32'h6f44e290, 32'h1309186, 32'h27c4d, 32'hb00009a, 32'h5a00c, 32'h0, 32'hb84e0, 32'h140302e0, 32'h0},{32'h0, 32'h0, 32'h8, 32'h1, 32'hc96c6000, 32'hcf366aa8, 32'h120309b, 32'h0, 32'h28400000, 32'h108810c, 32'h8b120010, 32'h20490, 32'h34000920, 32'h2},{32'h8000000, 32'h0, 32'hc00000, 32'h0, 32'h17b00000, 32'hb67a9422, 32'ha004ad, 32'h14003000, 32'h3000079, 32'h8611c, 32'ha000c000, 32'h18018000, 32'h7b0, 32'h0},{32'h2800, 32'h4040, 32'h0, 32'h0, 32'hc74ee2d0, 32'he19b7c8b, 32'h80a00145, 32'h27409, 32'h14c00004, 32'ha1008, 32'h8c000000, 32'h4000000, 32'h100108e0, 32'h0},{32'h0, 32'h0, 32'h1008, 32'h0, 32'h600003d0, 32'hf1cb54d1, 32'h5f038e4, 32'h5804800, 32'h23800078, 32'h213c, 32'h2f0c0000, 32'h1ec0f0, 32'h80000060, 32'h2},{32'h0, 32'h30, 32'h2000, 32'h0, 32'h15481618, 32'h23786bee, 32'h9e1393a, 32'h24802, 32'h1e400000, 32'h9e11c, 32'h9c0000a8, 32'h184020, 32'h0, 32'h0},{32'h0, 32'h20, 32'hca0000, 32'h4, 32'h94f4110, 32'hedb6ce20, 32'h5e02ce7, 32'h2384c, 32'h9447090, 32'h5e070, 32'h50, 32'h3a268000, 32'h740c0951, 32'h2},{32'h0, 32'h10, 32'h0, 32'h2, 32'h694f4000, 32'h2735662f, 32'h2001b8, 32'h0, 32'h2542908c, 32'h8c000, 32'h17000228, 32'h18228000, 32'h64020540, 32'h2},{32'h0, 32'h2000000, 32'h0, 32'h0, 32'h19686000, 32'hc249b2aa, 32'h8e000c5, 32'h11c27000, 32'h2504e095, 32'he000000, 32'h1c0a0184, 32'h0, 32'h680009c0, 32'h2},{32'h0, 32'h10030, 32'h2000, 32'h44000000, 32'h1d6c0e14, 32'h22aac51e, 32'h176, 32'h13c27800, 32'h12c4a094, 32'h4b000, 32'h0, 32'h74280, 32'h70000000, 32'h2},{32'h44, 32'h30, 32'h0, 32'h0, 32'h0, 32'h62adb000, 32'h9300b74, 32'h0, 32'h1c4e000, 32'h0, 32'h0, 32'h1e0000, 32'h70000910, 32'h2},{32'h0, 32'h40000000, 32'h4, 32'h0, 32'h0, 32'h72a81800, 32'h9713406, 32'h0, 32'h28000000, 32'ha0000, 32'h1f126000, 32'h170000, 32'h70000000, 32'h2},{32'h0, 32'h0, 32'hc02000, 32'h76000000, 32'hc18, 32'h50000000, 32'h212d24, 32'h0, 32'h12800000, 32'h7008, 32'h4a000000, 32'hf00bc000, 32'h600005d0, 32'h2},{32'h0, 32'h3004000, 32'h0, 32'h4, 32'h1470, 32'ha27a1000, 32'h92001b5, 32'h0, 32'h26800000, 32'h50089000, 32'h5c05c244, 32'h2824c170, 32'h341605c1, 32'h0},{32'h1000, 32'h0, 32'h4004, 32'h94000000, 32'hf6b, 32'hae341800, 32'h800001a4, 32'h3443, 32'h80600c, 32'h48090000, 32'h7114230, 32'h34450, 32'h30000000, 32'h0},{32'h8800000, 32'h0, 32'h0, 32'h0, 32'h68502000, 32'h49a87d51, 32'h2400114, 32'hf223400, 32'h5, 32'h0, 32'h0, 32'h180030, 32'h10000000, 32'h0},{32'h10000000, 32'h0, 32'h1000, 32'h0, 32'hc0000000, 32'h9a81e89, 32'h92054c2, 32'h13400000, 32'h2784d025, 32'h9c000, 32'h4000000, 32'h7c000, 32'h84010000, 32'h2},{32'h0, 32'h0, 32'h0, 32'h0, 32'ha546000, 32'h89c90cae, 32'h98001ad, 32'h13400000, 32'h1784f078, 32'h0, 32'h0, 32'hf42403d0, 32'h205003a0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h362041d0, 32'ha5766d14, 32'hc0015b, 32'h0, 32'h3000000, 32'h1a000, 32'h54124068, 32'h248060, 32'h64000000, 32'h0},{32'h4000000, 32'h280030, 32'h2010, 32'h0, 32'ha0000e10, 32'h71907d1b, 32'h98000c9, 32'h0, 32'h2340008d, 32'he800000, 32'h1d00022c, 32'h154000, 32'h0, 32'h0},{32'h11000, 32'h0, 32'h0, 32'h3, 32'hd0, 32'h0, 32'h80000000, 32'h2744a, 32'h86, 32'h88000, 32'h1c03c070, 32'h78000, 32'h442901e0, 32'h2},{32'h4000000, 32'h0, 32'h0, 32'h0, 32'hc0a78000, 32'h49507a9c, 32'h168, 32'h27c4e, 32'h26000095, 32'h0, 32'h240, 32'h228060, 32'h30000000, 32'h2},{32'h4000000, 32'h0, 32'h4280, 32'h0, 32'h1908, 32'hd18d4000, 32'h106, 32'h10c21800, 32'h9d, 32'h0, 32'h1c000000, 32'h1744e8, 32'h990, 32'h0},{32'h0, 32'h2, 32'h0, 32'h0, 32'h0, 32'h60000000, 32'h40a177, 32'h12825050, 32'h28425804, 32'ha0000, 32'h0, 32'h1704e0, 32'h20000880, 32'h2},{32'h0, 32'ha0000010, 32'h10, 32'h82000000, 32'ha000160e, 32'he6fbc218, 32'h126, 32'h0, 32'h1400000, 32'ha0000, 32'h2f0ba000, 32'h0, 32'h640009c0, 32'h2},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4000000, 32'h6000125, 32'h3000, 32'h60, 32'h8c000, 32'h5c000000, 32'h8000000, 32'h950, 32'h0},{32'h8000000, 32'h0, 32'h4, 32'h0, 32'h1810, 32'h6a4b1800, 32'h167, 32'hf000000, 32'hd, 32'h91000, 32'h8b05c180, 32'h0, 32'h984c0980, 32'h0},{32'h0, 32'h1000000, 32'h0, 32'h0, 32'h240, 32'haa0f0000, 32'h9b, 32'h13c00000, 32'h104e02c, 32'h0, 32'h1c, 32'h270000, 32'h9c0, 32'h0},{32'h0, 32'h0, 32'h4000, 32'h0, 32'h300001a0, 32'h72ac15d4, 32'hb, 32'h13c0e800, 32'h5e, 32'h0, 32'h7a0001e8, 32'h26c4e0, 32'h54000000, 32'h2},{32'hc000000, 32'h0, 32'h1010, 32'h2000000, 32'he0c, 32'haed0000, 32'h16c, 32'h1800000, 32'hb000091, 32'h0, 32'h55038070, 32'h1ec000, 32'h50000940, 32'h2},{32'h0, 32'h0, 32'h4, 32'h4, 32'h2b8, 32'h282fe060, 32'h8a, 32'h17000, 32'h5c, 32'h0, 32'h930a8000, 32'h0, 32'h6c000000, 32'h2},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'he0000000, 32'h167, 32'h0, 32'h0, 32'h0, 32'h5c000000, 32'h0, 32'h20000000, 32'h2},{32'h400c0, 32'h0, 32'h2000, 32'h0, 32'h110, 32'h0, 32'h9500087, 32'h27400, 32'h90, 32'h0, 32'h90010000, 32'h7c000, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h1, 32'h0, 32'hd8000000, 32'he7, 32'h0, 32'h26400000, 32'h0, 32'h0, 32'h0, 32'h34000000, 32'h2},{32'h10000140, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h500000, 32'h21c00, 32'h5, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h800, 32'h0, 32'h800000, 32'h0, 32'h0, 32'h0, 32'h80400000, 32'h1182844a, 32'h1846004, 32'h0, 32'h6000018, 32'h20000000, 32'h40000891, 32'h2},{32'h40000, 32'h0, 32'h0, 32'h0, 32'h475a0000, 32'h2eb6bbb5, 32'h41288b, 32'h1300344a, 32'h230290a1, 32'h0, 32'h0, 32'h0, 32'h40000000, 32'h2},{32'h0, 32'h0, 32'h10, 32'h0, 32'h10000000, 32'h5f35dd34, 32'h610008d, 32'h14027006, 32'h28000060, 32'h0, 32'h27114228, 32'h170000, 32'h0, 32'h0},{32'h40000, 32'h0, 32'h0, 32'h0, 32'h10000000, 32'hc298bd98, 32'hfc, 32'h1400, 32'h9c, 32'h8a000, 32'h200, 32'h0, 32'h990, 32'h0},{32'h80, 32'h5000000, 32'h10, 32'h0, 32'h1b0, 32'hf244e000, 32'h9f00102, 32'h1046, 32'h23000000, 32'h6000, 32'h7b00c1ec, 32'h25c000, 32'h0, 32'h0},{32'h8, 32'h0, 32'h0, 32'h1, 32'h0, 32'h65f89000, 32'h5f01b4c, 32'h0, 32'h26000000, 32'h8a000, 32'h7a0001e8, 32'h0, 32'h84460980, 32'h2},{32'h0, 32'h1008000, 32'h0, 32'h0, 32'hc0000000, 32'h52504a9d, 32'h5c100a8, 32'h0, 32'h0, 32'h40099000, 32'h7a00024c, 32'h0, 32'h950, 32'h0},{32'h0, 32'h0, 32'h10, 32'h0, 32'h1a00, 32'h6c000000, 32'h117, 32'h17400, 32'h0, 32'h0, 32'h1f05c000, 32'h258000, 32'h940, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'hb0000000, 32'ha7, 32'h1000, 32'h0, 32'h89130, 32'h1e000248, 32'h0, 32'h40000000, 32'h2},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4d180000, 32'h107, 32'h21800, 32'h0, 32'h88000, 32'h1e000000, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h48000000, 32'h9e00187, 32'h2784e, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'he8000000, 32'h18c, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h4000000, 32'h3000000, 32'h0, 32'h0, 32'h218, 32'h0, 32'h0, 32'h0, 32'h8d, 32'h0, 32'h5400001c, 32'h0, 32'h910, 32'h0},{32'h40, 32'h0, 32'h800000, 32'h0, 32'h0, 32'h70000000, 32'h950c017, 32'h0, 32'h99, 32'h0, 32'h0, 32'h0, 32'h8f0, 32'h0},{32'h4020100, 32'h0, 32'h0, 32'h0, 32'h1b10, 32'h0, 32'h9d00000, 32'h18400, 32'ha1, 32'h0, 32'h22c, 32'h0, 32'h0, 32'h0},{32'h0, 32'h10, 32'h0, 32'h0, 32'h0, 32'h0, 32'h9c00000, 32'h27850, 32'h22c50000, 32'h0, 32'h18, 32'h20c000, 32'h80000000, 32'h2},{32'h0, 32'h0, 32'h0, 32'h0, 32'h180, 32'h671a4000, 32'hc0015d, 32'h23400, 32'h0, 32'h90000, 32'h8a000000, 32'h0, 32'h0, 32'h0},{32'h100, 32'h0, 32'h2000, 32'h0, 32'h0, 32'h65a0000, 32'h5d000ed, 32'h0, 32'h0, 32'h0, 32'h0, 32'h264410, 32'h8000820, 32'h2},{32'h0, 32'h0, 32'h0, 32'h80d00000, 32'h802, 32'h0, 32'h8100000, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h5e0b800, 32'h17800, 32'h0, 32'h0, 32'h240, 32'h25c000, 32'hc0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'hea0a0800, 32'h18d, 32'h0, 32'h0, 32'h99000, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h89000, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h40, 32'h0, 32'h0, 32'h0, 32'h0, 32'h9f00000, 32'h0, 32'h1c00000, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h5c00000, 32'h13000000, 32'h180008c, 32'h0, 32'h0, 32'h20000000, 32'h8e1, 32'h0},{32'h100, 32'h0, 32'h0, 32'h0, 32'hc0000000, 32'h5ed45035, 32'h61000ba, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h5c000000, 32'h2},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h6000000, 32'h0, 32'h0, 32'h88130, 32'h0, 32'h258000, 32'h880, 32'h0},{32'h0, 32'h10000, 32'h0, 32'h0, 32'h0, 32'h4d5a9000, 32'hcd, 32'h0, 32'h0, 32'h7000, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h1, 32'h0, 32'h0, 32'h8400000, 32'h28400, 32'h22800000, 32'h0, 32'h0, 32'h0, 32'h84420000, 32'h2},{32'h0, 32'h10, 32'h1406000, 32'h4, 32'hca178000, 32'h7284e68d, 32'h93, 32'h23000, 32'h2640008c, 32'h6000, 32'h0, 32'h20c000, 32'hc468830, 32'h2},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h60000000, 32'h169, 32'h0, 32'h0, 32'h0, 32'h0, 32'h42104c0, 32'h10410841, 32'h2},{32'h0, 32'h0, 32'h0, 32'h0, 32'hc4254000, 32'hf1a9e216, 32'hd5, 32'h0, 32'h2284c000, 32'h6000, 32'h0, 32'h2084c0, 32'h80460900, 32'h1},{32'h0, 32'h0, 32'h0, 32'h0, 32'h10000800, 32'h568c4aa4, 32'h5f108d6, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4000000, 32'h18410861, 32'h2},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'hab694000, 32'h1b5, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h440000, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h99, 32'h0, 32'h0, 32'h2e000000, 32'h8f1, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h200, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h99112, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h4030000, 32'h0, 32'h8, 32'h0, 32'h0, 32'h0, 32'h0, 32'h22c00, 32'h8b, 32'h0, 32'h87000214, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h23400, 32'h0, 32'h0, 32'h84000210, 32'h0, 32'h960, 32'h0},{32'h0, 32'h0, 32'hc00004, 32'h87018004, 32'h21b, 32'h70000000, 32'ha2, 32'h3000, 32'h0, 32'h90000, 32'h99000264, 32'h0, 32'h84000850, 32'h1},{32'h0, 32'h0, 32'h0, 32'h1, 32'h0, 32'h8000000, 32'h12c, 32'h0, 32'h26400000, 32'h0, 32'h62000188, 32'h0, 32'h34300000, 32'h2},{32'h0, 32'h0, 32'h0, 32'h1, 32'h0, 32'hc0000000, 32'he4, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h1c000870, 32'h2},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h8a, 32'h0, 32'h88000000, 32'h0, 32'h18000000, 32'h2},{32'h0, 32'h6000000, 32'h4014, 32'h0, 32'hcb178000, 32'hf1c4e38d, 32'h82, 32'h0, 32'h0, 32'h0, 32'h85000214, 32'h214000, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h22800, 32'h2400008a, 32'h42000000, 32'h9710c050, 32'h210000, 32'h18000860, 32'h2},{32'h0, 32'h0, 32'h0, 32'h0, 32'haa400000, 32'h61117a18, 32'h166, 32'h0, 32'h1880008a, 32'h62110, 32'h88108210, 32'h0, 32'h30000000, 32'h2},{32'h0, 32'h0, 32'h0, 32'h0, 32'h1205, 32'h21cf9800, 32'h168, 32'h0, 32'h0, 32'h4c098000, 32'h9810818c, 32'h210000, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'hc9cc8800, 32'he7, 32'h0, 32'h26000000, 32'h0, 32'h98000210, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h50000000, 32'he8, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'hc0, 32'h1000020, 32'h0, 32'h0, 32'h0, 32'h0, 32'h8b00000, 32'h0, 32'h22400000, 32'h0, 32'h224, 32'h21c000, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h84000, 32'h0, 32'h0, 32'h78000000, 32'h2},{32'hc000000, 32'h10050, 32'h4, 32'h0, 32'hc0000000, 32'ha45e209, 32'h122, 32'h22c00, 32'h18c00091, 32'h63000, 32'h87000000, 32'h0, 32'h0, 32'h0},{32'h0, 32'h4000, 32'h0, 32'h0, 32'h0, 32'h0, 32'h9e00000, 32'h0, 32'h18800000, 32'h890c4, 32'h96000000, 32'h0, 32'h344f09a0, 32'h2},{32'h0, 32'h0, 32'h0, 32'h0, 32'h10000000, 32'h2934d3a6, 32'hea, 32'h0, 32'h0, 32'h99000, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h26400000, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h86000000, 32'h218000, 32'h0, 32'h0},{32'h0, 32'h0, 32'h40000, 32'h80100000, 32'hc03, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h3e000000, 32'h871, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h40, 32'h2000000, 32'h0, 32'h0, 32'h0, 32'h0, 32'h9f00000, 32'h0, 32'h0, 32'h0, 32'h264, 32'h0, 32'h9b0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h22800, 32'h0, 32'h0, 32'h220, 32'h0, 32'h9e0, 32'h0},{32'h0, 32'h6000000, 32'h4014, 32'h0, 32'hc5178000, 32'h7144e60d, 32'h103, 32'h0, 32'h0, 32'h0, 32'h8700021c, 32'h21c000, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h8a00000, 32'h22800, 32'h22000000, 32'h88000, 32'h86000220, 32'h218000, 32'h30000000, 32'h2},{32'h0, 32'h0, 32'h0, 32'h0, 32'h48324000, 32'h230cd41d, 32'h9e00187, 32'h0, 32'h26000000, 32'h43098000, 32'h86000260, 32'h34218000, 32'h9e1, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h48324000, 32'had51d41d, 32'h108, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h110c, 32'h0, 32'h0, 32'h0, 32'h0, 32'h22400, 32'h0, 32'h0, 32'h9f000000, 32'h27c468, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h22000, 32'h88, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h40, 32'hc000, 32'h0, 32'h87818000, 32'h21d, 32'h0, 32'h8b00000, 32'h0, 32'h0, 32'h89000, 32'h0, 32'h0, 32'h34000000, 32'h2},{32'h40, 32'hc020, 32'h0, 32'h0, 32'h0, 32'h0, 32'h9f00000, 32'h0, 32'h26400000, 32'h99000, 32'h0, 32'h0, 32'h9b0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h8a11800, 32'h0, 32'h0, 32'h0, 32'h0, 32'h278000, 32'h0, 32'h0},{32'h14060000, 32'h40, 32'h0, 32'h0, 32'hc6178000, 32'hf364e6cd, 32'h1a2, 32'h22400, 32'h22400089, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h8a11800, 32'h22000, 32'h22000088, 32'h0, 32'h9e000000, 32'h2304f0, 32'h300008e0, 32'h2},{32'h0, 32'h0, 32'h0, 32'h0, 32'hcd510000, 32'h29b476b0, 32'h9e001bb, 32'h11022000, 32'h26044098, 32'h98000, 32'h0, 32'h278000, 32'h9a0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'ha9568000, 32'h2a57b331, 32'h12c, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h3000000, 32'h2000, 32'h1, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h27c, 32'h23c000, 32'h3c0008d0, 32'h2},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h8c0, 32'h0},{32'h0, 32'h0, 32'h4, 32'h86000003, 32'ha18, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h9f000000, 32'h0, 32'h340008f0, 32'h2},{32'h4000080, 32'h30, 32'h0, 32'h0, 32'h0, 32'h0, 32'h9f00000, 32'h0, 32'h26400099, 32'h0, 32'h0, 32'h0, 32'h9b0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h1005000, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h234000, 32'h8d0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h9e00000, 32'h0, 32'h0, 32'h0, 32'h9e000278, 32'h18238460, 32'h380008e1, 32'h2},{32'h0, 32'h0, 32'h0, 32'h0, 32'hc42d4000, 32'he9cb821a, 32'he6, 32'h0, 32'h26000098, 32'h0, 32'h0, 32'h34230000, 32'h8c1, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h2e8ab000, 32'h146, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h1000000, 32'hc00000, 32'h0, 32'h218, 32'h0, 32'h9f00000, 32'h0, 32'h0, 32'h0, 32'h27c, 32'h0, 32'h8f0, 32'h0},{32'h4000000, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h99, 32'h0, 32'h0, 32'h0, 32'h9b0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h4000, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h23c000, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h9e00000, 32'h0, 32'h98, 32'h0, 32'h278, 32'h238000, 32'h9a0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h2a0cd000, 32'h166, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h9800000, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h80000000, 32'h2},{32'h40, 32'h0, 32'h0, 32'h34000000, 32'h808, 32'h0, 32'h9f00000, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h1400000, 32'h4, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h840009b0, 32'h2},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h28000, 32'ha0, 32'h0, 32'h0, 32'h0, 32'h80000000, 32'h2},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h60000000, 32'h164, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h28400, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h1, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0}};

