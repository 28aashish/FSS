//Constant array to load the A matrix
localparam integer A_size = 11;
localparam integer A[0:10] = '{32'h40a00000, 32'h40000000, 32'h3f800000, 32'h40800000, 32'hc0400000, 32'hc0a00000, 32'hc0000000, 32'hc0800000, 32'hbf800000, 32'h40c00000, 32'h40400000};
localparam integer A_BRAMInd[0:10] = '{0, 1, 2, 3, 0, 1, 0, 1, 2, 3, 2};
localparam integer A_BRAMAddr[0:10] = '{0, 0, 0, 0, 1, 1, 2, 2, 2, 2, 3};

//Constant array to load the instruction BRAM
localparam integer total_instructions = 56;
localparam integer sub_instructions = 10;
localparam integer Inst[0:55][0:9] = '{{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h200},{32'h0, 32'h0, 32'h22080000, 32'hc, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h80000000, 32'h4, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h40, 32'h0, 32'h20000000, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h40000, 32'h40000000, 32'h0, 32'h0},{32'h0, 32'h3000020, 32'h0, 32'h7480e80, 32'h2, 32'h0, 32'h10000, 32'h10000000, 32'h0, 32'h0},{32'h0, 32'h0, 32'h2000, 32'h4c00000, 32'h2, 32'h0, 32'h0, 32'h0, 32'h0, 32'h300},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h40, 32'h0, 32'h20000000, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h19443280, 32'h4, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h400},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h1000, 32'h4, 32'h0, 32'h0, 32'h30000, 32'h0, 32'h0, 32'h700},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h50000, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h20000, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h60000000, 32'h1, 32'h0, 32'h0, 32'h0, 32'h70000000, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h60000, 32'h0, 32'h0, 32'h600},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h2000, 32'h4c00000, 32'h1, 32'h0, 32'h0, 32'h0, 32'h0, 32'h500},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h20000, 32'h0, 32'h0, 32'h0, 32'h0, 32'h30, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h20, 32'h0, 32'h60000000, 32'h0, 32'h600},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h20800000, 32'h1, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h70000, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h70000000, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h1, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0}};

