//Constant array to load the A matrix
localparam integer A_size = 665;
localparam integer A[0:664] = '{32'h3e088c61, 32'hbd8888b5, 32'hb76ae18b, 32'hbd8888b5, 32'h3e088c61, 32'hbd8888b5, 32'hb76ae18b, 32'hbd8888b5, 32'h3e088ace, 32'hbd8888b5, 32'hbd8888b5, 32'hb70637bd, 32'h4170021b, 32'hb9fa9c13, 32'hb58637bd, 32'hb796feb5, 32'hb796feb5, 32'hb9fb224b, 32'h3b272eae, 32'hb8b88ca4, 32'hba828c37, 32'hba81a155, 32'hbd8888b5, 32'hbd8888b5, 32'h360637bd, 32'h390b75ea, 32'h3eaad2fe, 32'hb9712c28, 32'hbe4ccccd, 32'hb95f58c1, 32'hb76ae18b, 32'hb78637bd, 32'hbab02928, 32'h39ad8a11, 32'h3c51dcd7, 32'hbc441dd2, 32'h3955e8d5, 32'h3e08900c, 32'hbd8888b5, 32'hb7f34507, 32'hbd8888b5, 32'h3e088bdb, 32'hbd8888b5, 32'hbd8888b5, 32'hb75a1a93, 32'h40f00560, 32'hba19e0e7, 32'hb58637bd, 32'hb816feb5, 32'hb80a697b, 32'hba1aaa3b, 32'h3b81450f, 32'hba2d46f6, 32'hbad6909b, 32'hba8a8b09, 32'hbd8888b5, 32'hbd8888b5, 32'h368637bd, 32'h3948472c, 32'h3eaae4d2, 32'hb9d23d4f, 32'hbe4ccccd, 32'hb9798fa3, 32'hb7f34507, 32'hb81f6230, 32'hbb6874c9, 32'h3966afcd, 32'h3cd55821, 32'hbcc41dd2, 32'h3aa91538, 32'h3e088c61, 32'hb76ae18b, 32'hbd8888b5, 32'h3e088ace, 32'hbd8888b5, 32'hb716feb5, 32'h3cf3c2db, 32'hb87fda40, 32'hb58637bd, 32'hbcf2c301, 32'hb87fda40, 32'hb76ae18b, 32'hb8a5accd, 32'h3c69680e, 32'h3851b717, 32'hb78e9b39, 32'hbb113a50, 32'hbd8888b5, 32'hbd8888b5, 32'h36c9539c, 32'hb76ae18b, 32'h3eaaad1d, 32'h358637bd, 32'hb749539c, 32'hbcf2c301, 32'hb796feb5, 32'h3f5cedc4, 32'hb796feb5, 32'hbf555550, 32'h3d13165d, 32'hbcc41dd2, 32'hbc441dd2, 32'h3e08900c, 32'hbd8888b5, 32'hbd8888b5, 32'hb7f34507, 32'h3f800000, 32'hbd8888b5, 32'h3e088bdb, 32'hbd8888b5, 32'hb75a1a93, 32'hbd8888b5, 32'hbe4ccccd, 32'hbd8888b5, 32'h3eaaaf14, 32'hb6a7c5ac, 32'hb80a697b, 32'h36a7c5ac, 32'hb7f34507, 32'hbcc41dd2, 32'h358637bd, 32'h3cc4d445, 32'hb58637bd, 32'hb80e9b39, 32'hb7c9539c, 32'hb80637bd, 32'hb79f6230, 32'h3b8c2614, 32'hbb8b08dd, 32'h378e9b39, 32'hb80e9b39, 32'hbb8b08dd, 32'h3ed78983, 32'hb7e27e0f, 32'hbed55561, 32'hbcc41dd2, 32'hb75a1a93, 32'hb60637bd, 32'hb7e27e0f, 32'h3cc475e6, 32'hb716feb5, 32'hb851b717, 32'hbb0e25c8, 32'hb88e9b39, 32'hb7a7c5ac, 32'hbc441dd2, 32'h3c6a0ba2, 32'h3f800000, 32'h3e088c61, 32'hb76ae18b, 32'hbd8888b5, 32'hb76ae18b, 32'h3c449fd8, 32'hb78637bd, 32'h3e088a48, 32'hbd8888b5, 32'hb6c9539c, 32'h3bd6c2f0, 32'hb716feb5, 32'hb727c5ac, 32'hbbd6238e, 32'hbd8888b5, 32'hbd8888b5, 32'hb79f6230, 32'h3eaaad1d, 32'hb6c9539c, 32'hb727c5ac, 32'h3c449ba6, 32'hb76ae18b, 32'hbc441dd2, 32'hbf555550, 32'hb78637bd, 32'hbbd6238e, 32'hb76ae18b, 32'h3f57038e, 32'h40055554, 32'hbf555550, 32'h3f800000, 32'hbed55561, 32'hbf555550, 32'hbd8888b5, 32'h3e08900c, 32'hbd8888b5, 32'hb7f34507, 32'hbd8888b5, 32'h3e088d2a, 32'hbd8888b5, 32'hb796feb5, 32'hbe4ccccd, 32'hbd8888b5, 32'hbd8888b5, 32'h3eaaaf79, 32'hb7da1a93, 32'h377ba882, 32'hb7da1a93, 32'hbcc41dd2, 32'hb7f34507, 32'h38e27e0f, 32'h3ccfd8f1, 32'hb910b418, 32'hbaaf5fd4, 32'hb812ccf7, 32'hb6c9539c, 32'hb8e8c8ac, 32'h3c8f861a, 32'hb8e8c8ac, 32'hbc8da7f4, 32'hb796feb5, 32'hb910b418, 32'hbaa15981, 32'hb8dc3372, 32'h3cd0a244, 32'hb816feb5, 32'hbcc41dd2, 32'hbed55561, 32'hb816feb5, 32'hbc8da7f4, 32'hb816feb5, 32'h3ede392e, 32'h3cc41dd2, 32'hbc441dd2, 32'hbc441dd2, 32'h3e088c61, 32'hb76ae18b, 32'hbd8888b5, 32'hbc441dd2, 32'hb76ae18b, 32'h3c449fd8, 32'hb78637bd, 32'h3e088a48, 32'hb6eae18b, 32'hbd8888b5, 32'h3bd66f0d, 32'hb60637bd, 32'hb78637bd, 32'hbbd5cfab, 32'hb6eae18b, 32'h3c447a18, 32'hb60637bd, 32'hb76ae18b, 32'hbc441dd2, 32'hbd8888b5, 32'hbd8888b5, 32'hb79f6230, 32'h3eaaad1d, 32'hbf555550, 32'hb78637bd, 32'hbbd5cfab, 32'hb76ae18b, 32'h3f5702f7, 32'h3e088c61, 32'hb76ae18b, 32'hbd8888b5, 32'h3e088ace, 32'hbd8888b5, 32'hb716feb5, 32'h3cf02c4d, 32'hb896feb5, 32'hb60637bd, 32'hbceef805, 32'hb8991794, 32'hb76ae18b, 32'hb8dc3372, 32'h3c698138, 32'h385a1a93, 32'hb77ba882, 32'hbb101d19, 32'hbd8888b5, 32'hbd8888b5, 32'h36c9539c, 32'hb77ba882, 32'h3eaaad1d, 32'h3649539c, 32'hb749539c, 32'h3e088c61, 32'hb76ae18b, 32'hbd8888b5, 32'hb76ae18b, 32'h3c449fd8, 32'hb78637bd, 32'h3e088a48, 32'hbd8888b5, 32'hb6c9539c, 32'h3bd6ba8c, 32'hb727c5ac, 32'hb716feb5, 32'hbbd6238e, 32'hbd8888b5, 32'hbd8888b5, 32'hb79f6230, 32'h3eaaad1d, 32'hb6c9539c, 32'hb716feb5, 32'h3c449774, 32'hb76ae18b, 32'hbc441dd2, 32'hb78637bd, 32'hbbd6238e, 32'hb76ae18b, 32'h3f57038e, 32'hbf555550, 32'h3f800000, 32'h3e088c61, 32'hb76ae18b, 32'hbd8888b5, 32'hb76ae18b, 32'h3c449fd8, 32'hb78637bd, 32'h3bd6a9c5, 32'hb79f6230, 32'hbbd60a63, 32'h3e088a48, 32'hbd8888b5, 32'hb6eae18b, 32'hbd8888b5, 32'hb79f6230, 32'hbd8888b5, 32'h3eaaad1d, 32'hb6eae18b, 32'h3c4471b4, 32'hbc441dd2, 32'hb76ae18b, 32'hbc441dd2, 32'h3cc41dd2, 32'hbc441dd2, 32'hbf555550, 32'hb78637bd, 32'hbbd60a63, 32'hb76ae18b, 32'h3f57035c, 32'hbf555550, 32'h40055554, 32'hbf555550, 32'h3f800000, 32'hbed55561, 32'hbd8888b5, 32'h3e08900c, 32'hbd8888b5, 32'hb7f34507, 32'hbd8888b5, 32'h3e088d2a, 32'hbd8888b5, 32'hb796feb5, 32'hbe4ccccd, 32'hbd8888b5, 32'hbd8888b5, 32'h3eaaaf79, 32'hb7f34507, 32'h377ba882, 32'hb7c0f020, 32'hbcc41dd2, 32'hb7f34507, 32'h38e06530, 32'h3ccfce74, 32'hb910b418, 32'hbaae9681, 32'hb812ccf7, 32'hb6c9539c, 32'hb8e6afcd, 32'h3c8f1b26, 32'hb8e8c8ac, 32'hbc8d3cff, 32'hb796feb5, 32'hb910b418, 32'hbaa04d12, 32'hb8da1a93, 32'h3cd08f65, 32'hb816feb5, 32'hbcc41dd2, 32'hbed55561, 32'hb816feb5, 32'hbc8d3cff, 32'hb816feb5, 32'h3ede327f, 32'hbc441dd2, 32'hbcc41dd2, 32'h3f5e86b6, 32'hbf555550, 32'h3e088b54, 32'hbd8888b5, 32'hb7388ca4, 32'h3e088a48, 32'hbd8888b5, 32'hb6eae18b, 32'hbd8888b5, 32'hbd8888b5, 32'h3eaaac11, 32'hb727c5ac, 32'hb727c5ac, 32'h3b73eccc, 32'hbb734507, 32'h358637bd, 32'hb58637bd, 32'hbb734507, 32'h3f564ae0, 32'hb78e9b39, 32'hb78e9b39, 32'hbf555550, 32'hb6eae18b, 32'hb78e9b39, 32'h3c44827b, 32'hbc441dd2, 32'hbc441dd2, 32'hb7388ca4, 32'hb78e9b39, 32'hb58637bd, 32'h3c449774, 32'hbceef805, 32'hb796feb5, 32'hbf555550, 32'h3f5ccf5b, 32'hb796feb5, 32'hbc441dd2, 32'hb716feb5, 32'hb849539c, 32'hbb0dc11e, 32'hb890b418, 32'hb7b88ca4, 32'h3c69fadb, 32'hbc441dd2, 32'hbcc41dd2, 32'hbf555550, 32'h3f5e86b6, 32'hbc441dd2, 32'h3f5b763e, 32'hbf555550, 32'hbc441dd2, 32'h3e088c61, 32'hb76ae18b, 32'hbd8888b5, 32'h3e088ace, 32'hbd8888b5, 32'hb716feb5, 32'h3cf03afb, 32'hb88205ff, 32'hb58637bd, 32'hbcef3d3a, 32'hb8734507, 32'hb76ae18b, 32'hb8a17b0f, 32'h3c689a89, 32'h384d8559, 32'hb78e9b39, 32'hbb0e1501, 32'hbd8888b5, 32'hbd8888b5, 32'h36c9539c, 32'hb80a697b, 32'h3eaaacfb, 32'h358637bd, 32'h36eae18b, 32'hbcef3d3a, 32'hb796feb5, 32'h3f5cd196, 32'hb796feb5, 32'hbf555550, 32'h3d13165d, 32'hbc441dd2, 32'hbcc41dd2, 32'h3e088c61, 32'hbd8888b5, 32'hb76ae18b, 32'h3e088a48, 32'hbd8888b5, 32'hb6c9539c, 32'hbd8888b5, 32'hbd8888b5, 32'h3eaaacfb, 32'hb796feb5, 32'hb76ae18b, 32'h3c44a83b, 32'hb78e9b39, 32'hb60637bd, 32'hb75a1a93, 32'hb58637bd, 32'h3bd7a56e, 32'hbbd70e6f, 32'hb68637bd, 32'hb78e9b39, 32'hbbd70e6f, 32'h3f570564, 32'hb76ae18b, 32'hbf555550, 32'hbc441dd2, 32'hb6c9539c, 32'hb6a7c5ac, 32'hb76ae18b, 32'h3c4486ad, 32'hbd8888b5, 32'h3e08900c, 32'hbd8888b5, 32'hb7f34507, 32'hbd8888b5, 32'h3e088d2a, 32'hbd8888b5, 32'hb796feb5, 32'hbe4ccccd, 32'hbd8888b5, 32'hbd8888b5, 32'h3eaaaf79, 32'hb7da1a93, 32'h377ba882, 32'hb7da1a93, 32'hbcc41dd2, 32'hb7f34507, 32'h38dc3372, 32'h3ccfe154, 32'hb90d8ec9, 32'hbaafe60c, 32'hb816feb5, 32'hb68637bd, 32'hb8e8c8ac, 32'h3c90752e, 32'hb8e8c8ac, 32'hbc8e9d52, 32'hbcc41dd2, 32'hb796feb5, 32'hb910b418, 32'hbaa1dfb9, 32'hb8dc3372, 32'h3cd0a88f, 32'hb816feb5, 32'hb816feb5, 32'hbc8e9d52, 32'hb816feb5, 32'h3ede4884, 32'hbed55561, 32'hbf555550, 32'hbed55561, 32'h3fa4a287, 32'hbc441dd2, 32'hbcc41dd2, 32'h3cc41dd2, 32'hbc441dd2, 32'hbc441dd2, 32'h3e088c61, 32'hbd8888b5, 32'hb76ae18b, 32'h3e088ace, 32'hbd8888b5, 32'hb716feb5, 32'h3ced373b, 32'hb58637bd, 32'hb8841ede, 32'hb87fda40, 32'hbcec3116, 32'hbd8888b5, 32'hbd8888b5, 32'h36c9539c, 32'h3eaaacfb, 32'hb80205ff, 32'h36a7c5ac, 32'h358637bd, 32'hbc441dd2, 32'hb76ae18b, 32'hb8a9de8b, 32'h384d8559, 32'h3c684ad8, 32'hbb0ca3e8, 32'hb78e9b39, 32'hbc441dd2, 32'hb716feb5, 32'hb855e8d5, 32'hb88a697b, 32'hbb08722a, 32'h3c689eba, 32'hb7a7c5ac, 32'hb716feb5, 32'hb851b717, 32'hbb09a027, 32'hb88a697b, 32'hb7a7c5ac, 32'hbc441dd2, 32'h3c68ea3a, 32'hbf555550, 32'hbcec3116, 32'hb796feb5, 32'hb796feb5, 32'h3f5cb934, 32'hbf555550, 32'hbed55561, 32'hbc441dd2, 32'hbf555550, 32'h4006df33, 32'hbc441dd2, 32'hb75a1a93, 32'hb80a697b, 32'hb649539c, 32'hb58637bd, 32'hb58637bd, 32'hbcc41dd2, 32'h3cc486ad, 32'hb70637bd, 32'hb7b88ca4, 32'hba61f7d7, 32'hba102de0, 32'h39dbad3a, 32'hbc441dd2, 32'h3c54e4c9, 32'hbd8888b5, 32'h3e088ace, 32'hb716feb5, 32'hbd8888b5, 32'hbd8888b5, 32'hbd8888b5, 32'hbd8888b5, 32'hbe4ccccd, 32'hbc441dd2, 32'hbd8888b5, 32'hbd8888b5, 32'hbe4ccccd, 32'hbcc41dd2, 32'hbd8888b5, 32'h401e86b6, 32'hbd8888b5, 32'hbe4ccccd, 32'hbcc41dd2, 32'hbd8888b5, 32'hbd8888b5, 32'hbe4ccccd, 32'hbcc41dd2, 32'hbd8888b5, 32'hbd8888b5, 32'hbe4ccccd, 32'hbcc41dd2, 32'hbd8888b5, 32'hbd8888b5, 32'hbe4ccccd, 32'hbcc41dd2, 32'hbd8888b5, 32'h3f800000, 32'hbc441dd2, 32'hbe4ccccd, 32'h4170022d, 32'hba017fc7, 32'hb796feb5, 32'hb796feb5, 32'hb58637bd, 32'hba01c2e3, 32'h3b28e2e3, 32'hba8333fd, 32'hba82adc5, 32'hb8ae1049, 32'hb76ae18b, 32'hbc441dd2, 32'hb78637bd, 32'hbaac3a86, 32'h3c518d26, 32'h393fe3b0, 32'h39b2c83f, 32'hbc441dd2, 32'hb716feb5, 32'hb7b88ca4, 32'hba6cb74e, 32'h39ea5b53, 32'h3c558c8f, 32'hba1741d1, 32'hbd8888b5, 32'hbe4ccccd, 32'hbd8888b5, 32'h360637bd, 32'h390d8ec9, 32'hb9755de6, 32'hb969d51b, 32'h3eaad491};
localparam integer A_BRAMInd[0:664] = '{0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 5, 6, 1, 2, 3, 4, 5, 6, 0, 2, 3, 4, 5, 6, 7, 1, 2, 3, 4, 5, 6, 7, 0, 1, 3, 4, 5, 0, 1, 2, 3, 4, 5, 6, 7, 1, 2, 4, 5, 6, 7, 0, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 2, 3, 4, 5, 6, 7, 0, 1, 2, 4, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 4, 5, 7, 3, 4, 5, 6, 0, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 1, 2, 3, 4, 5, 6, 7, 0, 1, 3, 4, 5, 0, 1, 2, 3, 4, 5, 6, 0, 1, 2, 4, 5, 6, 7, 0, 1, 3, 4, 5, 6, 7, 0, 1, 2, 4, 5, 6, 1, 3, 4, 5, 6, 7, 1, 2, 3, 4, 6, 0, 2, 3, 4, 5, 6, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 1, 4, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 1, 2, 5, 6, 0, 3, 4, 5, 0, 1, 3, 4, 5, 6, 2, 3, 4, 5, 6, 7, 1, 3, 5, 0, 2, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 4, 6, 0, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 3, 4, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 4, 5, 6, 7, 0, 1, 3, 4, 5, 6, 7, 0, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 3, 4, 5, 6, 7, 0, 1, 3, 5, 6, 7, 0, 1, 2, 5, 1, 2, 4, 5, 7, 3, 4, 7, 2, 5, 7, 1, 2, 3, 4, 5, 7, 4, 7, 0, 1, 2, 3, 5, 7, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 7, 0, 1, 2, 6, 7, 0, 1, 2, 3, 4, 5, 0, 1, 2, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 3, 4, 5, 6, 7, 0, 1, 2, 3, 4, 5, 6, 7, 0};
localparam integer A_BRAMAddr[0:664] = '{0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 5, 5, 5, 5, 5, 6, 6, 6, 6, 6, 6, 6, 6, 7, 7, 7, 7, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 10, 10, 10, 10, 10, 10, 10, 10, 11, 11, 11, 11, 11, 11, 11, 11, 12, 12, 12, 12, 12, 12, 12, 13, 13, 13, 13, 13, 13, 13, 13, 14, 14, 14, 14, 14, 14, 14, 14, 15, 15, 15, 15, 15, 15, 15, 15, 16, 16, 16, 16, 16, 16, 16, 16, 17, 17, 17, 17, 17, 18, 18, 18, 18, 18, 18, 19, 19, 19, 19, 19, 19, 19, 20, 20, 20, 20, 20, 20, 20, 21, 21, 21, 21, 21, 22, 22, 22, 22, 22, 22, 22, 22, 23, 23, 23, 23, 23, 23, 24, 24, 24, 24, 24, 24, 24, 25, 25, 25, 25, 25, 25, 25, 25, 26, 26, 26, 26, 26, 26, 26, 26, 27, 27, 27, 27, 27, 27, 27, 27, 28, 28, 28, 28, 28, 28, 28, 28, 29, 29, 29, 29, 29, 29, 29, 30, 30, 30, 30, 30, 30, 31, 31, 31, 31, 31, 31, 31, 31, 32, 32, 32, 32, 32, 32, 33, 33, 33, 33, 34, 34, 34, 34, 34, 34, 35, 35, 35, 35, 35, 35, 35, 35, 36, 36, 36, 36, 36, 36, 36, 36, 37, 37, 37, 37, 37, 37, 37, 37, 38, 38, 38, 38, 38, 38, 38, 39, 39, 39, 39, 39, 40, 40, 40, 40, 40, 40, 40, 41, 41, 41, 41, 41, 41, 41, 42, 42, 42, 42, 42, 42, 42, 43, 43, 43, 43, 43, 43, 44, 44, 44, 44, 44, 44, 45, 45, 45, 45, 45, 46, 46, 46, 46, 46, 46, 47, 47, 47, 47, 47, 47, 47, 48, 48, 48, 48, 48, 48, 48, 48, 49, 49, 49, 49, 49, 49, 49, 49, 50, 50, 50, 50, 50, 50, 50, 50, 51, 51, 51, 51, 51, 51, 51, 51, 52, 52, 52, 52, 53, 53, 53, 53, 53, 53, 53, 53, 54, 54, 54, 54, 54, 54, 55, 55, 55, 55, 55, 55, 55, 56, 56, 56, 56, 57, 57, 57, 57, 58, 58, 58, 58, 58, 58, 59, 59, 59, 59, 59, 59, 60, 60, 60, 61, 61, 61, 61, 62, 62, 62, 62, 62, 62, 62, 62, 63, 63, 63, 63, 63, 63, 63, 63, 64, 64, 64, 64, 64, 64, 64, 64, 65, 65, 65, 65, 65, 65, 65, 66, 66, 66, 66, 66, 66, 66, 66, 67, 67, 67, 67, 67, 68, 68, 68, 68, 68, 68, 68, 69, 69, 69, 69, 69, 69, 69, 69, 70, 70, 70, 70, 71, 71, 71, 71, 71, 71, 71, 71, 72, 72, 72, 72, 72, 72, 72, 72, 73, 73, 73, 73, 73, 73, 73, 73, 74, 74, 74, 74, 74, 74, 74, 75, 75, 75, 75, 75, 75, 75, 76, 76, 76, 76, 76, 76, 77, 77, 77, 77, 77, 77, 77, 77, 78, 78, 78, 78, 78, 78, 78, 78, 79, 79, 79, 79, 79, 79, 79, 79, 80, 80, 80, 80, 80, 80, 80, 81, 81, 81, 81, 81, 81, 82, 82, 82, 82, 83, 83, 83, 83, 83, 84, 84, 84, 85, 85, 85, 86, 86, 86, 86, 86, 86, 87, 87, 88, 88, 88, 88, 88, 88, 89, 89, 89, 89, 89, 89, 89, 90, 90, 90, 90, 90, 90, 90, 90, 91, 91, 91, 91, 92, 92, 92, 92, 92, 93, 93, 94, 94, 94, 94, 96, 96, 96, 96, 96, 96, 96, 97, 97, 97, 97, 97, 97, 97, 97, 98, 98, 98, 98, 98, 98, 98, 99, 99, 99, 99, 99, 100, 100, 100, 100, 100, 100, 100, 100, 101};

//Constant array to load the instruction BRAM
localparam integer total_instructions = 914;
localparam integer sub_instructions = 12;
localparam integer Inst[0:913][0:11] = '{{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h21000000, 32'h84000, 32'h84000210, 32'h210000, 32'h380008e0, 32'h2},{32'h0, 32'h0, 32'h93980000, 32'ha44194, 32'h0, 32'h0, 32'h23800084, 32'h8e108, 32'h238, 32'h238000, 32'h38000000, 32'h2},{32'h0, 32'h0, 32'h44a00000, 32'h1485a6c, 32'h0, 32'h10400000, 32'h1780005e, 32'h0, 32'h5e000000, 32'h178000, 32'h704209c0, 32'h2},{32'h0, 32'h0, 32'ha3980000, 32'h9ba916, 32'h0, 32'h0, 32'h18, 32'h35000000, 32'h9a0d4178, 32'h2682f0, 32'h1a0, 32'h0},{32'h0, 32'h0, 32'h62ac0000, 32'h117c1ae, 32'h0, 32'h10400000, 32'h2680007c, 32'h9a000, 32'h0, 32'h8000000, 32'hf83506a1, 32'h1},{32'h0, 32'h0, 32'h4a2c0000, 32'hbbd24a, 32'h0, 32'h0, 32'h681d000, 32'h1a074, 32'h0, 32'h2703e0, 32'h700007c0, 32'h2},{32'h0, 32'h0, 32'h93100000, 32'h159b554, 32'h0, 32'h7800000, 32'hf000018, 32'h18000000, 32'h30000268, 32'h684d0, 32'h0, 32'h0},{32'h0, 32'h0, 32'ha32c0000, 32'h11741b7, 32'h0, 32'h0, 32'h1480007c, 32'h52000, 32'h3a138000, 32'he8000, 32'h700007e0, 32'h2},{32'h0, 32'h0, 32'h62ac0000, 32'h1493d0e, 32'h0, 32'h7400000, 32'hf000030, 32'h3a000, 32'h7c000000, 32'h0, 32'hc81f07c0, 32'h0},{32'h0, 32'h0, 32'h922c0000, 32'he52697, 32'h0, 32'h13000000, 32'h52, 32'h52000, 32'h0, 32'h8c0f8230, 32'h680003e0, 32'h2},{32'h0, 32'h0, 32'h93140000, 32'hd5a2f6, 32'h0, 32'hf800000, 32'h9a, 32'h30134, 32'h30094128, 32'h1f8000, 32'h0, 32'h0},{32'h0, 32'h0, 32'h9c9c0000, 32'h107b2f6, 32'h0, 32'hf800000, 32'h17800054, 32'h0, 32'h440fc110, 32'h0, 32'h802b0000, 32'h1},{32'h0, 32'h0, 32'hb2280000, 32'hfbc1c9, 32'h0, 32'h0, 32'h54, 32'h6a0a8, 32'h6a07c150, 32'hac000000, 32'h3e0, 32'h0},{32'h0, 32'h0, 32'h549c0000, 32'h1382ecf, 32'h0, 32'h0, 32'h0, 32'h4e04a0f8, 32'h4a0981f0, 32'h130000, 32'h70000000, 32'h2},{32'h0, 32'h0, 32'h849c0000, 32'h1143d93, 32'h0, 32'h0, 32'h4026010, 32'h12098, 32'h46000048, 32'h0, 32'h460, 32'h0},{32'h0, 32'h0, 32'h54a00000, 32'h159da8e, 32'h0, 32'h0, 32'h98, 32'h26044000, 32'h440000f8, 32'h34130000, 32'h3e1, 32'h0},{32'h0, 32'h0, 32'h549c0000, 32'h1162ed0, 32'h0, 32'h9800000, 32'h480001a, 32'h1a098, 32'h48, 32'h1a8000, 32'ha8000000, 32'h1},{32'h0, 32'h0, 32'h93100000, 32'h179d216, 32'h0, 32'h0, 32'h1f000030, 32'h23046000, 32'h1f0, 32'h64000000, 32'h460, 32'h0},{32'h0, 32'h0, 32'h55200000, 32'hbb4951, 32'h0, 32'h0, 32'h4022044, 32'h13000000, 32'h260000e8, 32'he8000, 32'h48000000, 32'h0},{32'h0, 32'h0, 32'h74180000, 32'h16aa291, 32'h0, 32'h0, 32'h15000012, 32'h2a026098, 32'h26000048, 32'h0, 32'h38000000, 32'h1},{32'h0, 32'h0, 32'h75a00000, 32'h89d232, 32'h0, 32'h0, 32'ha000000, 32'h28000, 32'h28000048, 32'ha0090, 32'h50000120, 32'h0},{32'h0, 32'h0, 32'h93980000, 32'h883554, 32'h0, 32'h0, 32'h11005028, 32'ha050, 32'ha0, 32'ha0000, 32'h18000000, 32'h1},{32'h0, 32'h0, 32'h62280000, 32'h169d650, 32'h0, 32'h0, 32'h600000a, 32'h18014, 32'h12000060, 32'h0, 32'h120, 32'h0},{32'h0, 32'h0, 32'h9ca00000, 32'h1483956, 32'h0, 32'h0, 32'h800000, 32'h28004, 32'h8, 32'h28000, 32'ha80000a0, 32'h0},{32'h0, 32'h0, 32'h82240000, 32'h1483153, 32'h0, 32'h0, 32'h2000008, 32'ha010, 32'h0, 32'h0, 32'h300000c0, 32'h0},{32'h0, 32'h0, 32'h92240000, 32'h169d26a, 32'h0, 32'h0, 32'h30000002, 32'h10c0000, 32'h28, 32'h4000000, 32'h80000a0, 32'h0},{32'h0, 32'h0, 32'h8c140000, 32'hb45256, 32'h0, 32'h0, 32'hc0, 32'h1000180, 32'h0, 32'h0, 32'h10000000, 32'h0},{32'h0, 32'h0, 32'h8ca00000, 32'h169d208, 32'h0, 32'h0, 32'h0, 32'hc0000, 32'h2000000, 32'h0, 32'h8610c20, 32'h0},{32'h0, 32'h0, 32'h93900000, 32'h1682a49, 32'h0, 32'h0, 32'h0, 32'h8000, 32'ha164000, 32'h590, 32'h500a0, 32'h0},{32'h0, 32'h0, 32'h93100000, 32'hf6b949, 32'h0, 32'h0, 32'h0, 32'h0, 32'h2c8, 32'h8590, 32'h8000000, 32'h0},{32'h0, 32'h0, 32'h4b100000, 32'ha4c1ae, 32'h0, 32'h5c00000, 32'h17017018, 32'h5c000, 32'h0, 32'h0, 32'h68180000, 32'h0},{32'h0, 32'h0, 32'haa2c0000, 32'h14926b7, 32'h0, 32'h0, 32'h21800000, 32'h0, 32'h0, 32'h218000, 32'h18440000, 32'h2},{32'h60000, 32'h1c050, 32'h10, 32'h52000000, 32'h5c50f8a1, 32'h83b10, 32'h2140008a, 32'h46090000, 32'h85120214, 32'h20240000, 32'h400008f1, 32'h2},{32'h1c040140, 32'h6000000, 32'h0, 32'h62000000, 32'h67ac92b1, 32'h138b3b10, 32'h23c00085, 32'h3208f0c8, 32'h180, 32'h23c300, 32'h78000000, 32'h2},{32'h180, 32'h1c000, 32'h4014, 32'h0, 32'h5444d300, 32'hd4d3c2e, 32'h1b80005f, 32'h60000, 32'h5f0c4000, 32'hc4180000, 32'h143609d0, 32'h2},{32'h80000000, 32'h18042, 32'h1c, 32'h30000000, 32'h592cafa1, 32'h172258, 32'h1f8450a0, 32'h2f87e140, 32'h9b0001ac, 32'h250000, 32'h580001b0, 32'h2},{32'h50000, 32'hc0000000, 32'h7010, 32'h6c000000, 32'h4c308899, 32'h123d2a, 32'h26c4f09e, 32'h8013c, 32'h9a000000, 32'hd6200200, 32'hfc500850, 32'h1},{32'h43000, 32'h5380000, 32'h0, 32'h30000000, 32'h5954e969, 32'h137598, 32'hec0d800, 32'h2009c064, 32'h32000070, 32'h1f44e8, 32'h700009e0, 32'h0},{32'h80000180, 32'h7000042, 32'h0, 32'hb0000000, 32'h55389389, 32'hfc83c24, 32'h3d, 32'h4d87e000, 32'hc4, 32'h406c1e0, 32'hf02a0541, 32'h0},{32'h40000, 32'h14c00, 32'h1c, 32'hf0000000, 32'h7ba48a59, 32'h83364, 32'h14c4003e, 32'h3e000, 32'h9d076000, 32'h782004a0, 32'h100007f0, 32'h2},{32'h180, 32'h10000, 32'h5380, 32'h2a000000, 32'h6c48b661, 32'hd4616, 32'h1582103b, 32'h42000, 32'h7d0ec1d8, 32'h158520, 32'hfc198000, 32'h0},{32'h180, 32'h4380000, 32'h5000, 32'h20000000, 32'h7ab4b879, 32'h94c3524, 32'hc825053, 32'h7e000, 32'h32000000, 32'h11c1f8, 32'h6c4004e0, 32'h2},{32'h1c000180, 32'h5000040, 32'h0, 32'h30000000, 32'h4bc8a951, 32'hc0e3d2a, 32'h1180009b, 32'h310fc, 32'h6000012c, 32'h1fc000, 32'h20000581, 32'h1},{32'h0, 32'h10050, 32'h6380, 32'h16000000, 32'h5428d899, 32'he3de8, 32'h6a, 32'h56084, 32'h7f0b0114, 32'h0, 32'h5c308580, 32'h1},{32'h10e00000, 32'h18000, 32'h14, 32'hb0000000, 32'h5c28af99, 32'h14d63e24, 32'h1280009c, 32'h550d6, 32'h3f13c000, 32'ha0298000, 32'h40000570, 32'h1},{32'h18e00000, 32'h14040, 32'h0, 32'h2e000000, 32'h47a0ab61, 32'h2943e2c, 32'h12000046, 32'h7d096, 32'h4d028274, 32'h90058000, 32'h28000140, 32'h1},{32'h1c040140, 32'h18000, 32'h0, 32'h90000000, 32'h65dcaca1, 32'ha2bec, 32'h13400011, 32'h13080, 32'h4709c278, 32'h140000, 32'h40000000, 32'h1},{32'h1c000000, 32'h43, 32'h14, 32'h18000000, 32'h6c3c9841, 32'h102e26, 32'h1a80e000, 32'h1f8450e4, 32'h16000134, 32'h2c070000, 32'hc80009b0, 32'h1},{32'h5010c, 32'h7000000, 32'h0, 32'he6000000, 32'h6aacae41, 32'h3743e18, 32'h4c2404d, 32'ha4144, 32'h800000c8, 32'h1ac000, 32'hd04104a0, 32'h0},{32'h14070000, 32'h60, 32'h10, 32'h94000000, 32'h74ccf2a9, 32'h10221c, 32'h1f413026, 32'ha0470ec, 32'h11c, 32'h281d8000, 32'hf0000330, 32'h0},{32'h80000100, 32'h63, 32'h5000, 32'h26000000, 32'h58d4d661, 32'h83e16, 32'h9828045, 32'h1d814054, 32'h9c, 32'ha4050000, 32'h4c0002a0, 32'h0},{32'h180501c0, 32'h0, 32'h4000, 32'h16000000, 32'h7928d3a9, 32'h5943618, 32'h1540a013, 32'h27000, 32'h90, 32'h48050000, 32'h3c1602c0, 32'h1},{32'h60000, 32'h501c000, 32'h4000, 32'h60000000, 32'h4adcd859, 32'h5893a98, 32'ha43a076, 32'h48000, 32'h290540e8, 32'h4c250, 32'h540002e0, 32'h0},{32'h50100, 32'h60, 32'h7000, 32'h14000000, 32'h6c5616b9, 32'h123b5e, 32'h2c42029, 32'h6016000, 32'he0000a4, 32'h1c030000, 32'h1c0b0860, 32'h1},{32'h1c040184, 32'h14200, 32'h3000, 32'h9c000000, 32'h5930d159, 32'h10eaa812, 32'h642900b, 32'h19000, 32'h1310e0a8, 32'h80102b0, 32'h244808e0, 32'h2},{32'h18440000, 32'h5004030, 32'h7000, 32'h98000000, 32'ha040f859, 32'h18dae12, 32'hc0605e, 32'h7003122, 32'h910c0234, 32'h2c060, 32'hac3906a0, 32'h0},{32'h8050100, 32'h0, 32'h7098, 32'h22000000, 32'h6034d5b9, 32'h89561f, 32'h2435009, 32'h6518c, 32'hc2000318, 32'hd4018610, 32'h344f80d0, 32'h0},{32'h4050186, 32'h8070, 32'h10, 32'h66000000, 32'h4634ae81, 32'hdf5582e, 32'h30450003, 32'h3f06100c, 32'h6300002c, 32'h381f04e0, 32'h18510031, 32'h0},{32'h1c250100, 32'h0, 32'h6100, 32'ha6000000, 32'hc0556341, 32'h18d56a62, 32'h44f0c1, 32'h6300111a, 32'h310, 32'h88298000, 32'h144b89c1, 32'h0},{32'h4000100, 32'h1c600, 32'h6114, 32'hae000000, 32'ha02cd089, 32'h138c562a, 32'h3202a001, 32'h81080, 32'h3082158, 32'h902701f0, 32'hc508c31, 32'h3},{32'h8000000, 32'h7010a00, 32'h6000, 32'he8000000, 32'hc0cda359, 32'h1850ae2e, 32'he802000, 32'h3033188, 32'hb3016074, 32'h90004000, 32'h2c6503c1, 32'h0},{32'h40, 32'h47018650, 32'h10, 32'h92000000, 32'h68dcd359, 32'h38aa02b, 32'h2380007f, 32'h4a09411c, 32'h11062cc, 32'haa00c000, 32'h784b0010, 32'h0},{32'h41984, 32'h200, 32'h5380, 32'h0, 32'h395ce800, 32'h7f1a263, 32'h1744082f, 32'h1a054060, 32'h9507a158, 32'hd0640, 32'hc40d8c80, 32'h0},{32'h10000, 32'h8030, 32'h0, 32'h0, 32'h38c24000, 32'h38a5b59, 32'h10c4208a, 32'h2704e094, 32'ha50001dc, 32'h980780d0, 32'h384604e0, 32'h1},{32'h40, 32'h3000000, 32'h2000, 32'h30b08000, 32'h54aa728a, 32'h8d76b2d, 32'hcc4504b, 32'h2d05408c, 32'h54090230, 32'h13c230, 32'h4420540, 32'h2},{32'h0, 32'h2000000, 32'hc, 32'h42e50000, 32'h2c5530bb, 32'h10979be3, 32'h61, 32'h1809c064, 32'h9a0680c8, 32'hc1641a0, 32'h78190811, 32'h2},{32'h46, 32'h8000, 32'h0, 32'hf0000000, 32'h99c9c85d, 32'h86d8be0, 32'h14026057, 32'h80000, 32'h59038200, 32'h41b4410, 32'h703f01a1, 32'h0},{32'hc0, 32'h4000, 32'h8, 32'h9e000000, 32'h96c13242, 32'h14ae16, 32'h118000a7, 32'h12088, 32'h9f000120, 32'h2c050000, 32'h34000510, 32'h1},{32'h0, 32'h0, 32'h0, 32'hc6000000, 32'h30ae4284, 32'h120c9029, 32'h2000004c, 32'h7c000, 32'h80000138, 32'h24238000, 32'h480008e1, 32'h2},{32'h0, 32'h180000, 32'h1000, 32'h84000000, 32'hc5dd4885, 32'h78e952e, 32'hf84f014, 32'h3e000, 32'h9c140270, 32'h284288, 32'hc090a00, 32'h1},{32'hc010000, 32'h0, 32'h0, 32'h44000000, 32'he54af4b2, 32'h1583ea, 32'h745101c, 32'h4f073000, 32'h6d0fc200, 32'h34000000, 32'h804d01e0, 32'h2},{32'h0, 32'h0, 32'hc, 32'hc4000000, 32'hb541e1ab, 32'ha514a2c, 32'h484e09a, 32'h0, 32'h7608c000, 32'h500504f0, 32'hd42a04b0, 32'h0},{32'h80, 32'h0, 32'h0, 32'hc6b10000, 32'h66b28173, 32'h949be2b, 32'h681b027, 32'h3d06c, 32'h2a050208, 32'h40883f0, 32'h30190221, 32'h1},{32'h4000000, 32'h0, 32'hc, 32'hc48b8000, 32'h9aaa8c73, 32'h134b6c26, 32'h480007e, 32'h3f015140, 32'h7c0000a0, 32'h440b0120, 32'ha4160531, 32'h0},{32'h10000, 32'h0, 32'h2000, 32'h6000000, 32'heb260c6d, 32'h13bae2, 32'h5424028, 32'h46000, 32'h5e0000a8, 32'hc41d8310, 32'hbc2302d0, 32'h0},{32'h0, 32'h0, 32'hc, 32'h44000000, 32'h2042c162, 32'h144b736b, 32'h205100c, 32'h53000000, 32'h86000218, 32'h2c2984e0, 32'h503f02f0, 32'h0},{32'h0, 32'h20, 32'h0, 32'h6e04000, 32'h9bad01b5, 32'h74c6c6a, 32'h1d000040, 32'h4809006c, 32'h90074034, 32'h6421c200, 32'he0000380, 32'h2},{32'h80, 32'h1180000, 32'h8000000, 32'hece0c432, 32'hb551f86d, 32'hc085e26, 32'h1804702b, 32'h13060084, 32'h571780f8, 32'h54244028, 32'h302200e0, 32'h0},{32'h20000, 32'h10, 32'h8000000, 32'h720d037, 32'h1c4e0952, 32'h24fae17, 32'h3402026, 32'h59000048, 32'h6c18c184, 32'hd81b0120, 32'h20140730, 32'h3},{32'hc000000, 32'h8000, 32'h3800000, 32'h9b2c0c, 32'h79d64100, 32'hf8a1b, 32'h28037080, 32'h400c70d4, 32'hc3144270, 32'h1f8380, 32'hb4400800, 32'h1},{32'hc010080, 32'h0, 32'h0, 32'h90a820, 32'h36c59600, 32'h91483eb, 32'h1fc000a1, 32'h2200714c, 32'h9c000120, 32'h298230, 32'h8c3a0740, 32'h2},{32'h46, 32'h20, 32'h0, 32'h0, 32'hd5423700, 32'h18ec74d2, 32'h2880009f, 32'h5e0a20f8, 32'ha708c314, 32'h1c1f85e0, 32'h903a0a41, 32'h2},{32'h21800, 32'h0, 32'h4, 32'hd0000000, 32'hfc518a94, 32'h15cd5c52, 32'h10464804, 32'h5903c018, 32'h3c1900f0, 32'h8060, 32'h640609f0, 32'h1},{32'h8000000, 32'h0, 32'h0, 32'h46e04012, 32'h99d9817c, 32'h17661a, 32'h5809046, 32'h230c5104, 32'h7e000190, 32'hf4240, 32'h98300820, 32'h1},{32'h4000000, 32'h0, 32'h100, 32'h50000000, 32'he9da2d82, 32'h254ae14, 32'h5800016, 32'h95024, 32'h24000058, 32'h30090000, 32'h5c0f8160, 32'h2},{32'h20000, 32'h10, 32'h0, 32'hec000000, 32'h78326ea4, 32'h16d4bad5, 32'h15c2804c, 32'h18002000, 32'h4e0980d4, 32'hc324000, 32'h48030b80, 32'h1},{32'hc0, 32'h0, 32'h1000, 32'hc4000000, 32'h1556c873, 32'h4992ef, 32'h1580504f, 32'h60056164, 32'hc000010, 32'h7c060, 32'h342b0040, 32'h2},{32'h4000000, 32'h20, 32'h3000, 32'h68018000, 32'h7836ae92, 32'h16d37c55, 32'h2704d032, 32'h505b060, 32'hb4014234, 32'h2185c0, 32'h241a0ac0, 32'h1},{32'h4000000, 32'h0, 32'h8000000, 32'h44365829, 32'h1c5e6da5, 32'h10a7e1d, 32'h681100e, 32'h23033030, 32'h350201d0, 32'h70000, 32'h883a0000, 32'h0},{32'h8000000, 32'h1000000, 32'h0, 32'h6000000, 32'h18227565, 32'h896bbd3, 32'h502a051, 32'h56081090, 32'h168, 32'h20c050, 32'h202e0ac0, 32'h1},{32'h0, 32'h2000000, 32'h0, 32'h145000, 32'h54cee300, 32'hca6c61, 32'hc83b02c, 32'h23032004, 32'h150ec200, 32'h5c170, 32'ha80407e0, 32'h0},{32'h30000, 32'h0, 32'h2004, 32'h81490000, 32'h86be3582, 32'h18179a6c, 32'h13c6303e, 32'h14178, 32'h14000318, 32'h802f0470, 32'h4c200930, 32'h2},{32'h20000, 32'h600, 32'h12c40004, 32'h1275849, 32'hd9800000, 32'h10bd58, 32'hfc0c0b8, 32'h9e000, 32'ha102e268, 32'h34290000, 32'h88300a11, 32'h0},{32'h0, 32'h0, 32'h2004, 32'hc6000000, 32'h5c4a0062, 32'h18164e11, 32'h2d06409c, 32'h7408c, 32'h9c028320, 32'ha82d80d0, 32'hc3a01f0, 32'h2},{32'hc000000, 32'h0, 32'h0, 32'h820589e0, 32'hd62672b3, 32'h10bd68, 32'ha005000, 32'h77000, 32'h160000a8, 32'h20048070, 32'h580800e0, 32'h0},{32'h10000, 32'h2000000, 32'h10, 32'h6000000, 32'h56a18e85, 32'h1649aad5, 32'hdc3f004, 32'hac00c, 32'h1200420c, 32'h4808c560, 32'h980604d0, 32'h0},{32'h0, 32'h2010030, 32'h0, 32'h901a8000, 32'hf9b5325b, 32'h177e2c, 32'h585c01a, 32'h2f046000, 32'h550ec094, 32'h740b40c0, 32'h505b0a31, 32'h0},{32'h20000, 32'h80000, 32'h0, 32'h86000000, 32'h15d10d7c, 32'h49b62b, 32'hac50006, 32'h4000, 32'h9c160020, 32'h818c258, 32'h10580a20, 32'h0},{32'h8000040, 32'hc000, 32'h0, 32'h94000000, 32'h882d12ab, 32'h9c9bbec, 32'h2e0000a3, 32'h200170a0, 32'hf0bc29c, 32'ha4138000, 32'hf85d04c0, 32'h0},{32'h80, 32'h0, 32'h4, 32'h6000000, 32'ha5b1578a, 32'h1d47a66, 32'h9004075, 32'h18020, 32'h560a82e4, 32'h18040000, 32'h60080390, 32'h1},{32'h0, 32'h1000030, 32'h2000, 32'hd0000000, 32'h56525873, 32'h95cef, 32'h8050bd, 32'h63000000, 32'hac00803c, 32'h80ac560, 32'h14030c20, 32'h1},{32'h4000000, 32'h0, 32'h0, 32'h80000000, 32'h5726828a, 32'hba3db, 32'h2d0070c0, 32'h61025000, 32'he000028, 32'h34028610, 32'h38000b60, 32'h0},{32'h80, 32'h1000000, 32'h0, 32'hd4000000, 32'haa18ea2, 32'h1cdb451, 32'h12003081, 32'h2000, 32'ha3000040, 32'h101c4230, 32'hc0050b00, 32'h2},{32'h0, 32'h20000000, 32'h10, 32'h44000000, 32'h35a24aa3, 32'h174c2b, 32'h1000000, 32'ha711c, 32'hbc00c000, 32'hea000000, 32'h290, 32'h0},{32'h0, 32'h1000000, 32'h4188, 32'h0, 32'h30000000, 32'h14abdd, 32'h2060008, 32'h5a0b4190, 32'h320, 32'h841d45a0, 32'h34528a51, 32'h1},{32'h4000000, 32'h1, 32'h0, 32'hc6000000, 32'h69369182, 32'h1850acdb, 32'h2880002a, 32'h380d000, 32'hc40002c4, 32'h500a8000, 32'h205207e0, 32'h1},{32'h4000000, 32'h0, 32'h180, 32'h240000, 32'hbb514900, 32'h176b98, 32'h22060086, 32'h83110, 32'h220, 32'h310000, 32'h64338c40, 32'h0},{32'h800000c0, 32'h10450, 32'h0, 32'h68000000, 32'h49d8b881, 32'h124aab20, 32'h2484a017, 32'hb892128, 32'h8704a21c, 32'h248000, 32'h48000190, 32'h2},{32'h18600000, 32'h20010050, 32'h2000, 32'h6e000000, 32'h4a4c9591, 32'h82b24, 32'h3003062, 32'h3109109e, 32'h91010244, 32'h72188320, 32'h4c320071, 32'h1},{32'h90051980, 32'h8000, 32'h0, 32'h9b410000, 32'h58d889b1, 32'hdd5bbd8, 32'h1842b861, 32'h286109c, 32'hd13c304, 32'he4138000, 32'h300009e0, 32'h1},{32'h800, 32'h611c000, 32'h4194, 32'hf0a1bc60, 32'h5c2cb8b9, 32'h128c44ee, 32'h2b45f81a, 32'h4801c128, 32'h6d000070, 32'h441b45c8, 32'ha44f86d0, 32'h0},{32'h0, 32'h610, 32'h4014, 32'h101c860, 32'h61000000, 32'hc138dd7, 32'h2c80000a, 32'h43062000, 32'h1103a1d4, 32'h682b0310, 32'h4460811, 32'h2},{32'h0, 32'h0, 32'h1100, 32'h80000000, 32'h79263865, 32'h14aadb, 32'hb00e06c, 32'h6c0c0, 32'h620381b0, 32'hd8188360, 32'h74258280, 32'h1},{32'h21800, 32'h0, 32'h0, 32'h83578000, 32'h374172a2, 32'h10d06d99, 32'h1dc40874, 32'h0, 32'h4010c010, 32'h10000, 32'h24440000, 32'h0},{32'h18200000, 32'h10050, 32'h0, 32'h71060000, 32'h4c38d8b1, 32'hc577a6c, 32'h31c300a2, 32'h4103d17a, 32'h3d10c0f4, 32'hc8208000, 32'h30400800, 32'h2},{32'h40, 32'h0, 32'h2000, 32'h86000000, 32'h55a1f8b2, 32'h84c4c6f, 32'h19061023, 32'h390640c0, 32'hbb078108, 32'h841b0610, 32'h844f0721, 32'h2},{32'h8000000, 32'h1000000, 32'h0, 32'he8348000, 32'hc8c1f794, 32'hd5d54, 32'h32400000, 32'h5075120, 32'h901242b8, 32'h582dc150, 32'ha0490921, 32'h0},{32'h0, 32'h1008000, 32'h0, 32'h6000000, 32'h37a5ca6a, 32'hb8c13, 32'h0, 32'h92120, 32'h17018030, 32'h3c120, 32'h504a0110, 32'h0},{32'h4400000, 32'h10000, 32'h0, 32'h1078000, 32'h81800000, 32'h10d29a5a, 32'h18000bf, 32'h715a, 32'h49110220, 32'hd8040, 32'h281b0000, 32'h2},{32'h10000146, 32'h2000000, 32'h6004, 32'h58000000, 32'h47c08849, 32'hef4ab6e, 32'h33, 32'h8716e, 32'h400000f0, 32'h64020, 32'hd4210bb0, 32'h0},{32'h0, 32'h10, 32'hc, 32'h268000, 32'h0, 32'hbce8240, 32'hb8, 32'h46086100, 32'hb1000024, 32'h0, 32'h30410a31, 32'h2},{32'h50086, 32'h20000000, 32'h10, 32'h0, 32'h28dae000, 32'h8335a51, 32'h540004f, 32'h94120, 32'h6c0001b0, 32'ha6000000, 32'h58370490, 32'h2},{32'h40080, 32'h1000000, 32'h3000, 32'h0, 32'h34000000, 32'h8107265, 32'hcc20025, 32'h11000, 32'h40078000, 32'h443d0, 32'h64000000, 32'h1},{32'h10000140, 32'h2000200, 32'h619c, 32'hb0000000, 32'h7c34b869, 32'hc8e7dea, 32'h1800003f, 32'h150c8, 32'h515a000, 32'h1c000, 32'h4648410, 32'h1},{32'h10000, 32'h8000, 32'hc, 32'h0, 32'h0, 32'h15d3a5c0, 32'h3c01006, 32'h2103c000, 32'hf06c30c, 32'h42c0000, 32'hd81a0b70, 32'h0},{32'hc0, 32'h4000050, 32'h8, 32'hd8000000, 32'h2c5aa1ba, 32'h484be3, 32'hc80a049, 32'h8816018, 32'hc000054, 32'h6c1540b0, 32'h181b0b10, 32'h0},{32'h0, 32'h10, 32'h0, 32'h1370000, 32'h45a2e000, 32'hc0dac93, 32'h15800080, 32'h800c8, 32'hb40ac2f4, 32'h282a0, 32'h330000, 32'h2},{32'h200100, 32'h0, 32'h3000, 32'h4000000, 32'h8b3db473, 32'h1813ba64, 32'hc81a07f, 32'ha0c916a, 32'h3402c0d0, 32'h58000, 32'h2c1a0c40, 32'h3},{32'h40, 32'h0, 32'h2000, 32'hc0000000, 32'h9aba9055, 32'hfcc8bdc, 32'h2000002b, 32'h1e0800b4, 32'h820b4108, 32'h2082a0, 32'h94220000, 32'h2},{32'h4030000, 32'h0, 32'h8, 32'he8000000, 32'hd9b2ee95, 32'hfd08a5e, 32'h224000a2, 32'h61089028, 32'hc2000058, 32'h483140b0, 32'h90400891, 32'h2},{32'h110c0, 32'h0, 32'h0, 32'h1170000, 32'h95dae800, 32'h64d9c2c, 32'h24c4a893, 32'ha034104, 32'h34048090, 32'h7024c410, 32'he0190801, 32'h2},{32'h0, 32'h3000010, 32'h2000, 32'he4000000, 32'h18355375, 32'h84adf, 32'h13000048, 32'h27074000, 32'h909018c, 32'he81943a0, 32'h94250480, 32'h1},{32'h0, 32'h200c000, 32'h1000, 32'h0, 32'ha6d9498d, 32'ha0b7c96, 32'hd819036, 32'h500ec, 32'h710081d8, 32'h1cc020, 32'hc4260480, 32'h1},{32'h10000, 32'h0, 32'h0, 32'hf68000, 32'h9bd2b600, 32'hdd054e4, 32'h8c21095, 32'h48000000, 32'h5a0a82f0, 32'h1c0360, 32'h70000400, 32'h1},{32'h4000000, 32'h2000030, 32'h0, 32'h58000000, 32'hf45558bb, 32'h108e1c, 32'h18836048, 32'h310630e4, 32'h480d82b4, 32'he4234250, 32'hb50, 32'h0},{32'h8000000, 32'h3004000, 32'h15020000, 32'h1514420, 32'he6800000, 32'h2cb7cec, 32'hd800032, 32'h6d028, 32'h63000050, 32'h300bc440, 32'he00c0880, 32'h0},{32'h0, 32'h60000000, 32'h88, 32'ha03400, 32'h4d2c800, 32'he979aef, 32'h76, 32'h62078, 32'h62000000, 32'hee000000, 32'h243b8430, 32'h2},{32'hc000000, 32'h44000000, 32'h4, 32'h1270000, 32'h0, 32'h179d80, 32'h1081603e, 32'h5e0a5178, 32'hc212020c, 32'h1a124000, 32'hb8140651, 32'h0},{32'h30000, 32'h10, 32'h0, 32'h70000, 32'hf9d2c200, 32'h15d54a22, 32'h1941b0b0, 32'h49024028, 32'h240041cc, 32'h702b0490, 32'hd00000c0, 32'h0},{32'hc000000, 32'h0, 32'h10000008, 32'h80d10451, 32'h39550b62, 32'h2d77d9d, 32'h503b048, 32'h2b000, 32'h240001d8, 32'h941200c0, 32'h930, 32'h0},{32'h40000, 32'h0, 32'h0, 32'h2000000, 32'hcad98b75, 32'h57a360, 32'h3415006, 32'h2a000, 32'h1d0, 32'h120000, 32'h54440740, 32'h2},{32'h0, 32'h3014000, 32'h2010, 32'h1590520, 32'h70000000, 32'h54a642d, 32'h782001e, 32'h2a000, 32'h9f03c000, 32'h3c0dc110, 32'h2c2009f0, 32'h2},{32'h14000000, 32'h40, 32'h0, 32'h71790000, 32'h4b552069, 32'h140b2be8, 32'h1800009e, 32'h1d000, 32'ha013c074, 32'h0, 32'h805109e0, 32'h2},{32'h0, 32'h10, 32'h100, 32'h30000000, 32'ha4d94815, 32'h167bae, 32'h78000a0, 32'he06c03c, 32'ha213c234, 32'h800f0, 32'hc5d81e0, 32'h2},{32'h40000, 32'h0, 32'h1000, 32'h18090000, 32'h16a893a1, 32'h167b95, 32'h743d000, 32'h53040000, 32'h3e14c070, 32'h3c1e8110, 32'h5c000401, 32'h2},{32'h80000000, 32'h1008041, 32'h0, 32'haa000000, 32'hc49c062, 32'hf5c5b, 32'h780d0b4, 32'h3d81c164, 32'h7b000014, 32'h10c000, 32'h805b0b60, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h55524800, 32'h14d35d93, 32'h806065, 32'h60020, 32'ha613c000, 32'h20000000, 32'hc05d0ba0, 32'h2},{32'h0, 32'h44000000, 32'h4, 32'h6000000, 32'h2539f745, 32'hc0bacd3, 32'h880e0bc, 32'h90000, 32'h371742f0, 32'h1227c110, 32'he8000450, 32'h2},{32'h0, 32'h8000, 32'h4, 32'h0, 32'h2b36b400, 32'h13c8bbe1, 32'h56, 32'h5901714c, 32'h714c300, 32'h40278000, 32'h60600371, 32'h1},{32'h80020040, 32'h41, 32'h0, 32'h1612040, 32'hc9dd8b00, 32'h6898c1e, 32'h15c07081, 32'h5a816184, 32'h34, 32'h18308000, 32'h9c6100e0, 32'h1},{32'h0, 32'h620, 32'h0, 32'h115c52, 32'hba800000, 32'h140c4cd4, 32'h10800080, 32'h0, 32'h1718a0d4, 32'h278000, 32'h8200a20, 32'h2},{32'h10230000, 32'h8000, 32'h0, 32'h161a060, 32'h90000000, 32'h185762a8, 32'h2040000a, 32'h50b6, 32'h8302c000, 32'h40000, 32'h40620000, 32'h0},{32'h0, 32'h0, 32'h2004, 32'h78000, 32'h66000000, 32'h175251, 32'h32, 32'h6006008, 32'he0000d0, 32'hc038000, 32'h94000a50, 32'h2},{32'h8000000, 32'h10, 32'h0, 32'h380000, 32'h1702d800, 32'hb9c99, 32'h1380004e, 32'h2083164, 32'h1000c094, 32'hc300000, 32'h40060b90, 32'h0},{32'h600000, 32'h1000000, 32'h2000, 32'h141d860, 32'h17a12e00, 32'h136b17, 32'hc800000, 32'h607509e, 32'hac1642b0, 32'h1d45c0, 32'h2c600b80, 32'h1},{32'h44, 32'h0, 32'h0, 32'h0, 32'h182a8d00, 32'h6e97e1d, 32'h51, 32'h4077008, 32'h2e0, 32'h0, 32'hd0040b80, 32'h0},{32'h0, 32'h2180000, 32'h1000, 32'h0, 32'h88000000, 32'h99c54, 32'h2f400000, 32'h0, 32'hb0000010, 32'h114388, 32'h74250b00, 32'h1},{32'h10000000, 32'h0, 32'h0, 32'h148000, 32'h0, 32'ha8380, 32'hc6, 32'hd0e6, 32'hc6164000, 32'h0, 32'h700d01c0, 32'h0},{32'h0, 32'h0, 32'h1100, 32'h0, 32'hfb000000, 32'h84a9c, 32'h0, 32'h700c158, 32'h481581d8, 32'h38000, 32'h641c8190, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h28c1c000, 32'h190f94d9, 32'h2c80000c, 32'h1c, 32'hc8164000, 32'h0, 32'hd0050000, 32'h2},{32'h4000080, 32'h0, 32'h0, 32'h0, 32'h99d24800, 32'he7dec, 32'h3000043, 32'hbd188, 32'hac000000, 32'h84000000, 32'hbc000c41, 32'h0},{32'h4000000, 32'h40, 32'h8, 32'h0, 32'h41800000, 32'ha5cdd, 32'h900c0b1, 32'h25000, 32'h30c, 32'h0, 32'h28000390, 32'h1},{32'h10000, 32'h0, 32'h0, 32'h240000, 32'h0, 32'h14a8c0, 32'h1dc63000, 32'h610c6000, 32'hc4000010, 32'h64620, 32'h20000000, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h17220100, 32'h128d5b, 32'h320000b0, 32'h610c8000, 32'h1d4, 32'h0, 32'hc0020000, 32'h2},{32'h40, 32'h10030, 32'h2000, 32'h0, 32'h9b000000, 32'h128d10, 32'h1f, 32'h0, 32'h503e08c, 32'h280000, 32'hc000000, 32'h1},{32'h0, 32'h3000000, 32'h1100, 32'hc10040, 32'h0, 32'h0, 32'h19000066, 32'hf066000, 32'h1e0dc198, 32'hcc2ec370, 32'h8c5086e0, 32'h2},{32'h43980, 32'h1180050, 32'h8000000, 32'hd6e0c422, 32'h67c0b2a1, 32'h110a2354, 32'h1b43186d, 32'h88000, 32'ha311418c, 32'h7c108, 32'h8a0, 32'h0},{32'h30080, 32'h5004000, 32'h10, 32'h0, 32'h57800000, 32'hd922dd4, 32'h1ec33041, 32'h3301c000, 32'h2300829c, 32'h10224380, 32'hc0040890, 32'h1},{32'h10000000, 32'h0, 32'h2004, 32'hb0000000, 32'h76c4950c, 32'hc897ad1, 32'h188320b5, 32'h63000, 32'h40c8188, 32'h60000000, 32'h84320b71, 32'h0},{32'h40080, 32'h0, 32'h4, 32'h86000000, 32'hb86985b, 32'hd89a3eb, 32'h30c490a7, 32'h3901112c, 32'h96000258, 32'h281c8000, 32'hbb1, 32'h0},{32'h20040, 32'h4014060, 32'h0, 32'h66000000, 32'h65b89071, 32'hcbc6a, 32'h8c440bd, 32'h880c4, 32'h9317624c, 32'h1024c320, 32'h80320c01, 32'h2},{32'h4000000, 32'h0, 32'h0, 32'h240140, 32'hba800000, 32'h99b64, 32'h3049000, 32'ha7000, 32'hc2124228, 32'h10038450, 32'h500008a1, 32'h2},{32'h40000, 32'h14000, 32'h0, 32'h2070000, 32'hb6a8b065, 32'h157a14, 32'hac49092, 32'h490bc000, 32'h89058188, 32'hc8248000, 32'h900002c0, 32'h1},{32'h100, 32'h0, 32'h1000, 32'h1e000000, 32'h5d59651, 32'h12928e11, 32'h2504b02b, 32'h49088000, 32'h8812c030, 32'h20248000, 32'h14450a30, 32'h1},{32'h0, 32'h0, 32'h0, 32'h2000000, 32'hcbc9c95c, 32'h7cf8d68, 32'h25020040, 32'h0, 32'h8c1241b8, 32'h18220000, 32'h144b06e1, 32'h3},{32'h0, 32'h4400, 32'h4000, 32'h20000000, 32'hf4ad8e51, 32'h555bda8, 32'h18800066, 32'h7018, 32'hf172198, 32'h800b8000, 32'hbc170101, 32'h1},{32'h0, 32'h4000, 32'h0, 32'h58000, 32'h4b2a6200, 32'h9bb21, 32'h19000000, 32'h620e4, 32'h7110230, 32'h10230390, 32'h983708c1, 32'h1},{32'h0, 32'h2000010, 32'h0, 32'hd8000000, 32'h2429f052, 32'hd4ce9, 32'h25036000, 32'h49000000, 32'hc10e42b4, 32'he02e4390, 32'hc0000960, 32'h1},{32'h80000000, 32'h0, 32'h0, 32'h0, 32'h55d22a00, 32'hdabd1, 32'ha85e0bc, 32'h5c8bc000, 32'h70124024, 32'hb0490, 32'hc03702c0, 32'h1},{32'h0, 32'h0, 32'h0, 32'h5c000000, 32'hdaaa8c42, 32'h127da4, 32'h16815000, 32'h5a0b0, 32'hb1000070, 32'h6c1605b0, 32'hb80002e1, 32'h0},{32'h102, 32'h0, 32'h5000, 32'h66000000, 32'h55489461, 32'h18eb8351, 32'h57, 32'h38000, 32'he0000d8, 32'h6c2e0000, 32'h641d01d0, 32'h1},{32'h18040144, 32'h0, 32'h0, 32'h170000, 32'h54b0b800, 32'heeb2c24, 32'hd400035, 32'h3101715a, 32'ha008320, 32'hc2e8030, 32'h38610ba0, 32'h0},{32'h100, 32'h0, 32'h5100, 32'h40000000, 32'h1621c182, 32'hacb7b55, 32'h3081a081, 32'h0, 32'h5806c000, 32'h3102c0, 32'hc5a8360, 32'h2},{32'h80000000, 32'h40, 32'h0, 32'h0, 32'h77328000, 32'h6caabdb, 32'he01a080, 32'h57838104, 32'h8200005c, 32'h70000000, 32'h90410a40, 32'h2},{32'h10000000, 32'h0, 32'h0, 32'h28000000, 32'h99a2ca91, 32'h717aadc, 32'hd000080, 32'hb035070, 32'h50104208, 32'h30000000, 32'h9c0c0500, 32'h0},{32'h40140, 32'h2004000, 32'h0, 32'h5c000000, 32'h15bed051, 32'h6d3a5d3, 32'h13c6384f, 32'h4068, 32'hc5000000, 32'h6c0241b0, 32'he0000b00, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h36aa4100, 32'h9d79a17, 32'h32427050, 32'hb0a4048, 32'h90, 32'ha4140000, 32'h90410500, 32'h2},{32'h0, 32'h0, 32'h0, 32'h58000000, 32'h75a13255, 32'h108ced, 32'h1381a050, 32'h6e02c, 32'h2e0, 32'h605c0, 32'h480c0000, 32'h1},{32'h8000000, 32'h4000000, 32'hc, 32'h104800, 32'h365a8800, 32'hdac13, 32'h2c8000b4, 32'h670b4, 32'h0, 32'h12c378, 32'h702c0670, 32'h1},{32'h0, 32'h4000, 32'h0, 32'h0, 32'h94000000, 32'hed4bda6, 32'h89, 32'h740ec, 32'h8b000000, 32'h1d0250, 32'h0, 32'h0},{32'h20000, 32'h100c000, 32'h0, 32'h0, 32'hd9000000, 32'h6936dd8, 32'h19c00036, 32'h160c4, 32'hb7174090, 32'h741c41c0, 32'h98000091, 32'h0},{32'h40, 32'h3000020, 32'h0, 32'h0, 32'h245aed00, 32'h164b9be1, 32'h7000065, 32'h3416c, 32'h651702ec, 32'h42c45c0, 32'hd0000b60, 32'h2},{32'hc000000, 32'h1, 32'h4, 32'h0, 32'h49b64f00, 32'h175a15, 32'h30800088, 32'h4b89718c, 32'h1cc, 32'h0, 32'h20000950, 32'h3},{32'h10000, 32'h0, 32'h10, 32'h1608000, 32'h0, 32'h13a200, 32'h22461000, 32'hc8000, 32'he000000, 32'h194000, 32'h280004b0, 32'h3},{32'h0, 32'h1000020, 32'h0, 32'h370000, 32'h0, 32'h12aa00, 32'h1d800000, 32'h76000, 32'h6400022c, 32'h9422c320, 32'h54000940, 32'h2},{32'h80, 32'hc000, 32'h8000004, 32'ha1342e, 32'h0, 32'h125d00, 32'h22000093, 32'h3a000000, 32'h2d148298, 32'h941d0000, 32'hfc510650, 32'h2},{32'h40, 32'h4194000, 32'h0, 32'h302a0000, 32'h4c3cb881, 32'h3cc5c52, 32'h25c10095, 32'h20000, 32'ha1040080, 32'h84284088, 32'h8000200, 32'h1},{32'h98000000, 32'h10451, 32'h1000, 32'haa802c00, 32'h483cb279, 32'h12572a9e, 32'h41, 32'h3781f000, 32'h1f11a07c, 32'h0, 32'h5c4a0000, 32'h2},{32'h40, 32'h8000, 32'h0, 32'h9b8000, 32'h0, 32'h3c00000, 32'h67, 32'h0, 32'h1103c1b8, 32'hbc370, 32'h80000000, 32'h0},{32'h0, 32'h3000020, 32'h1000, 32'h1068000, 32'h0, 32'h177a00, 32'h8800040, 32'h1107303c, 32'h2203c234, 32'h234210, 32'h9c000000, 32'h1},{32'h0, 32'h40000000, 32'h4, 32'hdb0000, 32'hf8800000, 32'he9d1c, 32'h1e, 32'h1e000, 32'h730580b0, 32'h2e080000, 32'h711, 32'h0},{32'h10000, 32'h200c000, 32'h0, 32'hf14040, 32'h0, 32'h169300, 32'h2f4000bd, 32'h0, 32'h71148078, 32'hb4000, 32'h0, 32'h0},{32'hc020000, 32'h20000050, 32'h10, 32'h0, 32'hc000000, 32'hf2601, 32'h16c000a6, 32'h53059000, 32'ha2140304, 32'h5e2dc000, 32'h88000a10, 32'h2},{32'h10400000, 32'h0, 32'h1000, 32'h0, 32'hf7000000, 32'h117d90, 32'h0, 32'h30c3172, 32'h601c0dc, 32'h40000000, 32'hec510a21, 32'h0},{32'hc0, 32'h80000, 32'h0, 32'he009f1, 32'h0, 32'h95a80, 32'hc9, 32'h5305814c, 32'hc4000160, 32'h1c5d8, 32'ha00, 32'h0},{32'h0, 32'h200, 32'h70000000, 32'h100c822, 32'h0, 32'h1154c0, 32'h0, 32'h6184, 32'h370b2310, 32'h18620, 32'h0, 32'h0},{32'h4030000, 32'h40000000, 32'h0, 32'h1260000, 32'h0, 32'hd9c00, 32'he441000, 32'h83044, 32'h18044078, 32'h4a000000, 32'h391, 32'h0},{32'h0, 32'h400c020, 32'h4, 32'h1513820, 32'h0, 32'h18cf84c0, 32'h39, 32'h1b0c6184, 32'h5106c20c, 32'h304000, 32'h190, 32'h0},{32'h80, 32'h1000000, 32'h0, 32'hf0c420, 32'h0, 32'h129dc0, 32'hb1, 32'h41082000, 32'ha40a0140, 32'hdc500, 32'he4000000, 32'h0},{32'h0, 32'h3000000, 32'h18000004, 32'h128bc70, 32'h0, 32'he6880, 32'h0, 32'h25000, 32'hb603c000, 32'h301445b0, 32'h530, 32'h0},{32'h0, 32'h0, 32'h2000, 32'h158000, 32'h0, 32'h190d7b80, 32'hb2, 32'hc8184, 32'h2e4, 32'h8000, 32'h4c000000, 32'h1},{32'h0, 32'h0, 32'h1000, 32'h0, 32'hc0000000, 32'h129dec, 32'h0, 32'h0, 32'h0, 32'h0, 32'h74000000, 32'h1},{32'h4000000, 32'h40, 32'h0, 32'h0, 32'h0, 32'h0, 32'h77, 32'h75000, 32'h3c, 32'h0, 32'h0, 32'h0},{32'h0, 32'h2000000, 32'h1000, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'hbb020038, 32'he4080, 32'h9c000000, 32'h0},{32'h4000000, 32'h8000, 32'h0, 32'h0, 32'h0, 32'hd83c0, 32'h0, 32'h70b7158, 32'hb90002b0, 32'h0, 32'hd4000000, 32'h2},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h108cc0, 32'h0, 32'hb603c, 32'h0, 32'h2d8000, 32'h24000000, 32'h3},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'hc9c80, 32'h0, 32'h70b4000, 32'h2d0, 32'h0, 32'h2c000000, 32'h3},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h108c80, 32'h1dc00000, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h21800, 32'h1000000, 32'h0, 32'h0, 32'h0, 32'h0, 32'h29453800, 32'h78000, 32'h720001d4, 32'h28c000, 32'he8000700, 32'h1},{32'h14430000, 32'h10010, 32'h0, 32'h50000000, 32'h5c38b891, 32'h122614, 32'h8400000, 32'h6f042, 32'h6f000084, 32'h0, 32'h210, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h6e0e41c8, 32'he01c0000, 32'h200, 32'h0},{32'h0, 32'h0, 32'h0, 32'ha00000, 32'he6000000, 32'hf7416, 32'h0, 32'h0, 32'h0, 32'h0, 32'h84000000, 32'h0},{32'h0, 32'h10, 32'h0, 32'h0, 32'h0, 32'h0, 32'h8c00000, 32'h0, 32'h8c, 32'h0, 32'h80000000, 32'h0},{32'h0, 32'h0, 32'h0, 32'h40000, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h80000100, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h89, 32'h5b800000, 32'h294, 32'h0, 32'h0, 32'h0},{32'h40000, 32'h4000, 32'h0, 32'h0, 32'h0, 32'h11000000, 32'h3c000a7, 32'h0, 32'ha3114000, 32'h228000, 32'h0, 32'h0},{32'h0, 32'h5018000, 32'h10, 32'h0, 32'h0, 32'hcbbc0, 32'h3800088, 32'h56000000, 32'h651182b8, 32'h46194460, 32'h951, 32'h0},{32'h0, 32'h0, 32'h4000, 32'h0, 32'h67800000, 32'hc91a41b, 32'h25800094, 32'ha7000, 32'h7a188258, 32'h28190000, 32'h2c330961, 32'h2},{32'h0, 32'h0, 32'h4014, 32'h70078000, 32'hba596a71, 32'hcd76260, 32'h64, 32'h46066000, 32'h64000228, 32'hcc228460, 32'hc450430, 32'h1},{32'h0, 32'h0, 32'h4000, 32'h60000000, 32'he5b53162, 32'h1275ec, 32'h42, 32'h230f0, 32'h7a1741e8, 32'h842e8320, 32'h54210440, 32'h2},{32'h0, 32'h40, 32'h0, 32'h30000000, 32'h98596a99, 32'hecc6bdc, 32'h198000c7, 32'h4b0960cc, 32'h1bc, 32'h190000, 32'hd84a0420, 32'h1},{32'h0, 32'h4000000, 32'h0, 32'h30000000, 32'hca453241, 32'h855e6, 32'h94, 32'ha50e4, 32'h720001b8, 32'hf010c000, 32'h584a02e0, 32'h2},{32'h0, 32'h10050, 32'h0, 32'h30000000, 32'h9428b859, 32'he84ec, 32'h2f0070bc, 32'h10000, 32'h2d16e0b4, 32'h2d0080, 32'h284a0000, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h9b310100, 32'h84daca8, 32'h1e8000c9, 32'h0, 32'h700f41b8, 32'h110210, 32'h10210700, 32'h1},{32'h0, 32'h0, 32'h0, 32'h50000000, 32'hd62a0eba, 32'hf6d2e, 32'h2f807000, 32'h5a000000, 32'h2c0c82e8, 32'h5c0b85d0, 32'hd8210760, 32'h1},{32'h14000000, 32'h10060, 32'h0, 32'h54000000, 32'hf82dcc42, 32'h11ad1a, 32'h1602d058, 32'hf000, 32'h700001c, 32'h0, 32'h0, 32'h0},{32'h14c00000, 32'h40, 32'h0, 32'h0, 32'h4c50b800, 32'h1425aa, 32'h2f000000, 32'h5918a, 32'h1100c164, 32'h10020000, 32'hf8000940, 32'h2},{32'h10000000, 32'h0, 32'h0, 32'h0, 32'ha4000000, 32'hb7b28, 32'h0, 32'h300715a, 32'hb000c2c0, 32'h682c0000, 32'hd0000a41, 32'h2},{32'h40000, 32'h14000, 32'h0, 32'h30000000, 32'hf5b1ee51, 32'hc8c10, 32'h20c2d000, 32'hb70b0, 32'h19010018, 32'h0, 32'h70000080, 32'h1},{32'h0, 32'h10050, 32'h0, 32'h0, 32'h34000000, 32'ha83eb, 32'h1a000000, 32'hb5000, 32'h370000dc, 32'h2a8000, 32'h48000680, 32'h1},{32'h10000000, 32'h14060, 32'h0, 32'h30000000, 32'h5c28d461, 32'h17c83614, 32'hb0, 32'h1608300c, 32'h51150144, 32'h2c0000, 32'hd0000780, 32'h2},{32'h1000, 32'h4000010, 32'h0, 32'h30000000, 32'h3b2a2379, 32'h89dd9, 32'h1e439800, 32'h1b0a4104, 32'h360001c4, 32'h700641c0, 32'he0000a40, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'he5aa7200, 32'h88b50, 32'he000038, 32'h1b070000, 32'h5006c1c0, 32'h0, 32'h481d0520, 32'h1},{32'h0, 32'h1000000, 32'h0, 32'h100c820, 32'hfb21ca00, 32'h148a68, 32'h0, 32'h24154, 32'h181501cc, 32'h1c40c0, 32'h98000000, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'hec49a800, 32'hf74e4, 32'h31864000, 32'h1b0b8188, 32'hb806c2e0, 32'h0, 32'h20650000, 32'h3},{32'h0, 32'h0, 32'h0, 32'he0000000, 32'h343a3273, 32'h159a69, 32'h0, 32'h800601c, 32'h20, 32'h40000, 32'h80, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h28000000, 32'hc9c55, 32'h2b000000, 32'he000, 32'h2b0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h109500, 32'h0, 32'h8a000, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h1200000, 32'h0, 32'h0, 32'h0, 32'h0, 32'h8b000000, 32'h0, 32'h0, 32'h0},{32'h0, 32'h4000, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h8d0002bc, 32'h198000, 32'h0, 32'h0},{32'hc010000, 32'h0, 32'h8, 32'hc00000, 32'h0, 32'h0, 32'h25c00000, 32'h7b000, 32'h8a000000, 32'h0, 32'h9c000970, 32'h1},{32'h0, 32'h20, 32'h4, 32'h370000, 32'h0, 32'h0, 32'h67, 32'h0, 32'h234, 32'h0, 32'h670, 32'h0},{32'hc0, 32'h40000010, 32'h10, 32'h0, 32'h0, 32'h0, 32'h79, 32'h0, 32'hbb0001ec, 32'h8a000000, 32'h210, 32'h0},{32'h8010000, 32'h0, 32'h3000, 32'h0, 32'h0, 32'h0, 32'h19c00077, 32'h5b097040, 32'hb6000080, 32'hcc000000, 32'he4330200, 32'h1},{32'h0, 32'h4188000, 32'h1000, 32'hb48000, 32'ha9800000, 32'he5460, 32'h0, 32'h11073044, 32'h2f020018, 32'h843c8, 32'h5c5a0200, 32'h2},{32'h40, 32'h0, 32'h0, 32'h78000, 32'h1000000, 32'h1154d3, 32'h80110bd, 32'h110b6000, 32'hb6000080, 32'h1c0100, 32'h440, 32'h0},{32'h0, 32'h0, 32'h18003000, 32'h262861, 32'hdac1b400, 32'he6ca2, 32'h1ec00000, 32'h0, 32'h2e000000, 32'h0, 32'h14000000, 32'h1},{32'h0, 32'h2000010, 32'hc, 32'he10000, 32'h0, 32'h0, 32'h2fc00000, 32'h0, 32'h2ec, 32'hb40bc000, 32'h770, 32'h0},{32'h2, 32'h0, 32'h0, 32'h202c00, 32'h0, 32'hb600000, 32'h59, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h40, 32'h1000, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h314, 32'h24000, 32'hfc000000, 32'h2},{32'hc0, 32'h8000, 32'h4, 32'h0, 32'h0, 32'h18c00000, 32'h318000a5, 32'h62000000, 32'hb10002c4, 32'h20000, 32'hb50, 32'h0},{32'h0, 32'h0, 32'h1000, 32'h60000, 32'h0, 32'h148dc0, 32'h320000c8, 32'h0, 32'h310, 32'h0, 32'h74000000, 32'h1},{32'h20000, 32'h1000600, 32'h0, 32'h0, 32'h0, 32'h148580, 32'h1a400000, 32'h0, 32'h53156000, 32'h1a4000, 32'h0, 32'h0},{32'h30002, 32'h0, 32'h2000, 32'h0, 32'h0, 32'h16200000, 32'h2a4000bf, 32'h0, 32'h38000000, 32'h0, 32'hec000000, 32'h1},{32'h8000000, 32'h0, 32'h4, 32'hb820, 32'h0, 32'h0, 32'h0, 32'ha5000, 32'h52000000, 32'h148000, 32'h390, 32'h0},{32'h40, 32'h0, 32'h8, 32'he13040, 32'h0, 32'h0, 32'h20800039, 32'h0, 32'h0, 32'h2a8000, 32'hec000530, 32'h0},{32'h0, 32'h0, 32'h2004, 32'h0, 32'h0, 32'hca000, 32'h0, 32'h0, 32'h0, 32'h0, 32'h9c000270, 32'h0},{32'h8000000, 32'h30, 32'h80, 32'h0, 32'h0, 32'h0, 32'h0, 32'hb9000, 32'h100002e4, 32'h20000, 32'h2c648000, 32'h3},{32'h0, 32'h0, 32'h0, 32'h1601c0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h2b400000, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h1e0000a8, 32'h0, 32'h1c8, 32'h0, 32'h0, 32'h0},{32'h14000000, 32'h40, 32'h0, 32'h0, 32'h5c589800, 32'h102e28, 32'h0, 32'h71000, 32'h1c4, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h1c83c020, 32'h38000000, 32'h1c8, 32'h0, 32'he8000000, 32'h1},{32'h4000000, 32'h0, 32'h0, 32'h1608000, 32'h1a000000, 32'h158a21, 32'h0, 32'h21000, 32'hb40142dc, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'he7840, 32'h0, 32'h23040, 32'h0, 32'h0, 32'h0, 32'h0},{32'h10000, 32'h0, 32'h0, 32'h298000, 32'h0, 32'h0, 32'h8c00000, 32'hb7000, 32'h8c000260, 32'h0, 32'h60000000, 32'h2},{32'h10000000, 32'h0, 32'h0, 32'h0, 32'h48000000, 32'he2610, 32'h0, 32'h8b000, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h19800000, 32'h0, 32'hba000000, 32'h0, 32'h0, 32'h0},{32'h0, 32'h4000000, 32'h0, 32'h0, 32'h4c000000, 32'h14261c, 32'h0, 32'h0, 32'h0, 32'h19c000, 32'h60000000, 32'h2},{32'h0, 32'h40, 32'h0, 32'h0, 32'h0, 32'h82600, 32'h1a000000, 32'h34000000, 32'h22c, 32'h198000, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h116500, 32'hc7, 32'h45000000, 32'h8c000230, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'he8c00, 32'hc9, 32'h0, 32'h1a0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h10, 32'h0, 32'h0, 32'h102600, 32'h0, 32'h0, 32'h0, 32'h0, 32'h670, 32'h0},{32'h10000000, 32'h0, 32'h0, 32'h0, 32'h0, 32'hcc00000, 32'h198000a8, 32'h11000, 32'hba0002e8, 32'h0, 32'h660, 32'h0},{32'h0, 32'h6010000, 32'h14, 32'h0, 32'habd89800, 32'he5428, 32'ha8, 32'h7005c, 32'h71000000, 32'h114000, 32'h450, 32'h0},{32'h0, 32'h10000, 32'h0, 32'h0, 32'h4c000000, 32'hed69026, 32'h1c00005a, 32'h72000, 32'h2f0e01c8, 32'h88000000, 32'h760, 32'h0},{32'h0, 32'h0, 32'h4014, 32'h30000000, 32'h5958b8a1, 32'ha5de8, 32'h1e83c078, 32'h570ac020, 32'h700001e8, 32'hec110000, 32'h6c3c05b0, 32'h1},{32'h0, 32'h0, 32'h0, 32'h12000000, 32'heb41945b, 32'h129c6a, 32'h5a, 32'h7a000, 32'h1e8, 32'h0, 32'h702d0440, 32'h1},{32'h0, 32'h0, 32'h0, 32'h0, 32'h94000000, 32'h1054ac, 32'h2f800000, 32'hb4020, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h10000, 32'h0, 32'h0, 32'h0, 32'h129d00, 32'h0, 32'h0, 32'h9000000, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'hb00102c0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'he7c00, 32'h38, 32'h0, 32'h780002e0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h4014000, 32'h0, 32'h0, 32'h4c40b800, 32'h162e1c, 32'h0, 32'h0, 32'h390b8000, 32'he42e0, 32'h0, 32'h0},{32'h0, 32'h45010000, 32'h4, 32'h0, 32'h57800000, 32'h70d261a, 32'h73, 32'hb8000, 32'h530002e0, 32'h5614c1c0, 32'he80007b1, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'hd4000000, 32'h106cae, 32'h0, 32'h0, 32'h2e000000, 32'h1e0000, 32'h0, 32'h0},{32'h10000, 32'h0, 32'h0, 32'h0, 32'h0, 32'hc7000, 32'h1cc00000, 32'h0, 32'h8000000, 32'h1a0290, 32'hb40, 32'h0},{32'h80000000, 32'h42, 32'h0, 32'h0, 32'he0000000, 32'hc6e14, 32'h0, 32'h8800000, 32'h24, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h17c00000, 32'h2b0000b0, 32'h80ac000, 32'hb0000020, 32'h0, 32'hb40, 32'h0},{32'h0, 32'h10, 32'h0, 32'h0, 32'hbba1600, 32'h128d15, 32'h23400000, 32'h0, 32'h264, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h4000000, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'hbb000, 32'h0, 32'h0, 32'ha4000000, 32'h1},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h52000000, 32'h1a0000, 32'h990, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'hc7000, 32'h23000000, 32'h8c000, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h1205000, 32'h0, 32'h0, 32'h0, 32'h5b022000, 32'h234, 32'h0, 32'h0, 32'h0},{32'h100, 32'h0, 32'h0, 32'h0, 32'h4c000000, 32'h122622, 32'h21, 32'h69000, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h2a0, 32'h0, 32'ha0000000, 32'h1},{32'h40040, 32'h0, 32'h2000, 32'h808000, 32'h0, 32'h4102600, 32'h8417067, 32'h54000000, 32'h2ec, 32'h0, 32'hac000000, 32'h2},{32'h0, 32'h0, 32'h0, 32'h1a8000, 32'h0, 32'h11b800, 32'h8810000, 32'h5b02216c, 32'h700001c8, 32'h0, 32'h0, 32'h0},{32'h6, 32'h0, 32'h8, 32'h0, 32'h5a41c100, 32'he31ace5, 32'h77, 32'h0, 32'h0, 32'h0, 32'h5d0, 32'h0},{32'h20040, 32'h0, 32'h3000, 32'h0, 32'h0, 32'h0, 32'h1ec00079, 32'h0, 32'h2bc, 32'h0, 32'he40005c0, 32'h1},{32'h0, 32'h0, 32'h1000, 32'ha08000, 32'h0, 32'h0, 32'h0, 32'h7b000, 32'h0, 32'h0, 32'h74000000, 32'h1},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h2fc00000, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h2c4, 32'h0, 32'h0, 32'h0},{32'h0, 32'h10, 32'h2000, 32'h0, 32'h0, 32'h0, 32'h0, 32'h5c000, 32'h1e4, 32'h0, 32'hf40003b0, 32'h2},{32'h0, 32'h4000, 32'h0, 32'h90000, 32'h0, 32'h0, 32'h0, 32'h0, 32'h5d000000, 32'h0, 32'h3a0, 32'h0},{32'h0, 32'h0, 32'h1000, 32'ha08000, 32'h0, 32'h0, 32'h0, 32'hb9000, 32'h78070000, 32'h0, 32'hec000000, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'he7800, 32'h0, 32'he000, 32'h2d0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h109040, 32'h0, 32'h0, 32'h69000000, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h44, 32'h0, 32'h0, 32'h0, 32'h0, 32'h16200000, 32'h2b4000bf, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h1a400000, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h4000000, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'hbf000, 32'h0, 32'h0, 32'h94000000, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'ha9000, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h22, 32'hab000, 32'h0, 32'h0, 32'h90000000, 32'h0},{32'h410000, 32'h0, 32'h0, 32'h160a020, 32'h0, 32'h0, 32'h8c00000, 32'hb70e6, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h94000000, 32'h0, 32'h980, 32'h0},{32'h10050000, 32'h0, 32'h0, 32'h0, 32'h4c000000, 32'he2e14, 32'h23400000, 32'h8d000, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h23000000, 32'h8c000, 32'h94000260, 32'h0, 32'h58000980, 32'h2},{32'h0, 32'h0, 32'h0, 32'h0, 32'h24000000, 32'haa41d, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h4000, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'ha4000000, 32'h1},{32'h0, 32'h0, 32'h10, 32'h0, 32'h0, 32'h0, 32'h1a000000, 32'h68174, 32'h2e8, 32'h0, 32'ha0000310, 32'h1},{32'h0, 32'h0, 32'h0, 32'h0, 32'h8a000000, 32'h1044e4, 32'h0, 32'hb4000, 32'h40, 32'h0, 32'hec000000, 32'h1},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h128000, 32'h0, 32'h0, 32'h170, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h10, 32'h0, 32'h0, 32'h102600, 32'h0, 32'h0, 32'h0, 32'h0, 32'h5d0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h70, 32'h72000, 32'h0, 32'h0, 32'h5c0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h165480, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h100, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h5d, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h10, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h3b0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'hb8000, 32'h1e0, 32'h0, 32'he85e03a0, 32'h1},{32'h0, 32'h0, 32'h0, 32'h0, 32'ha4000000, 32'h125260, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h80000, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h25c4c8, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h258000, 32'h960, 32'h0},{32'h0, 32'h0, 32'h1000, 32'ha0b020, 32'h0, 32'h0, 32'h0, 32'h0, 32'h264, 32'h0, 32'h5c000000, 32'h2},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h68, 32'hb6000, 32'h0, 32'h0, 32'h0, 32'h0},{32'h10100, 32'h0, 32'h5000, 32'h1608000, 32'h0, 32'h122600, 32'h1a45a023, 32'hbb000, 32'h0, 32'h0, 32'h940d0000, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h4554800, 32'h2a000024, 32'h5c150, 32'h0, 32'h0, 32'h98120260, 32'h0},{32'h0, 32'h0, 32'h0, 32'h90000, 32'h955ae800, 32'h13bd2c, 32'h0, 32'haa150, 32'h0, 32'h0, 32'h90000000, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h134480, 32'h1c800072, 32'hbe16c, 32'h0, 32'h0, 32'h90000000, 32'h0},{32'h0, 32'h0, 32'h0, 32'h1405800, 32'h0, 32'h134480, 32'h0, 32'h73000, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h80, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'hf43d8000, 32'h2},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h2dc00000, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'hb5, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h2000, 32'h110000, 32'h0, 32'h0, 32'h2a400000, 32'h0, 32'h0, 32'h0, 32'h9c000000, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'hab000, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'hbf000, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h17800000, 32'h96, 32'h96000, 32'h98000000, 32'h260000, 32'h0, 32'h0},{32'h0, 32'h5000000, 32'h10, 32'h0, 32'h475cb800, 32'h122d98, 32'h0, 32'h0, 32'h0, 32'h25c000, 32'h970, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h258000bc, 32'h96000, 32'h260, 32'h2604b0, 32'hf8000960, 32'h2},{32'h0, 32'h0, 32'h0, 32'h0, 32'hd8495400, 32'h165218, 32'h0, 32'hba000, 32'h0, 32'h0, 32'h0, 32'h0},{32'h100, 32'h0, 32'h0, 32'h0, 32'h0, 32'h122600, 32'h69, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h68, 32'h0, 32'h740001d0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h4000, 32'h0, 32'h0, 32'heb400, 32'h0, 32'h0, 32'h0, 32'h0, 32'h7c000000, 32'h1},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h40140, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h1cc00073, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'he400000, 32'h1c800078, 32'haa000, 32'h0, 32'h54000000, 32'he85507a1, 32'h1},{32'h0, 32'h0, 32'h0, 32'h10000000, 32'h45daeab5, 32'h9bc93, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h4000, 32'h8, 32'h0, 32'h0, 32'h0, 32'h97, 32'h0, 32'h99000000, 32'h0, 32'hbf0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h96, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h20000, 32'h10, 32'h0, 32'h1610000, 32'h0, 32'h0, 32'h25c00000, 32'h0, 32'h264, 32'h0, 32'hfc000000, 32'h2},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h2ec00000, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h74000, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h10, 32'h1200000, 32'h0, 32'h0, 32'h0, 32'h0, 32'h1d4, 32'h0, 32'h270, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h2d800000, 32'hbe000, 32'h0, 32'h0, 32'h260, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h145480, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h2a000000, 32'h0, 32'h0, 32'h0, 32'h260, 32'h0},{32'h0, 32'h0, 32'h3004, 32'h218000, 32'h0, 32'h145000, 32'h0, 32'h0, 32'h0, 32'h0, 32'hec000ab0, 32'h1},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'hbf000, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'hab000, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h100, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h97, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h96, 32'h0, 32'h98000260, 32'h0, 32'hf8000be0, 32'h2},{32'h0, 32'h0, 32'h0, 32'h0, 32'h68000000, 32'h8b29d, 32'h2e800000, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h10000000, 32'h0, 32'h0, 32'h0, 32'h0, 32'h142600, 32'h0, 32'h75000, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h1d800076, 32'h74000, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h149580, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h10, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h7b0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'haa17c, 32'h0, 32'hf4000000, 32'hf0000aa0, 32'h2},{32'h0, 32'h0, 32'h0, 32'h0, 32'hb9000000, 32'h85cd4, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h26000000, 32'h98000, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h10, 32'h0, 32'h120d020, 32'h0, 32'h0, 32'h0, 32'h0, 32'h264, 32'h0, 32'hbf0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'hbb, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'he0000000, 32'h1},{32'h0, 32'h0, 32'h0, 32'h800000, 32'h0, 32'h0, 32'h77, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h200000, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'hbf156, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'hac, 32'h0, 32'h280, 32'h0, 32'hbe0, 32'h0},{32'h10050000, 32'h0, 32'h0, 32'h0, 32'h4c289800, 32'h102e2c, 32'h26400000, 32'h99000, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h2605f0ac, 32'h57098000, 32'h280, 32'h7c000000, 32'ha21, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h48c24a00, 32'hba56d, 32'hba, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h4000, 32'h0, 32'h0, 32'h162600, 32'h0, 32'h0, 32'h0, 32'h0, 32'he4000000, 32'h1},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h1e800000, 32'h7a000, 32'h0, 32'h0, 32'he0000000, 32'h1},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h124500, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h2000000, 32'h1000, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h28c, 32'h2fc000, 32'hbc000000, 32'h2},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'ha2000288, 32'h288000, 32'h0, 32'h0},{32'h0, 32'h10, 32'h10000008, 32'hc13850, 32'h0, 32'h0, 32'h2fc00000, 32'h0, 32'h2bc, 32'h0, 32'ha30, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'hbd0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h7a, 32'h0, 32'h0, 32'h0, 32'hf0000000, 32'h1},{32'h0, 32'h0, 32'h0, 32'h1602000, 32'h0, 32'h0, 32'h1ec00000, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'ha6000, 32'h290, 32'h0, 32'hb8000000, 32'h2},{32'h0, 32'h4014060, 32'h0, 32'h70000000, 32'h4c48d841, 32'h103610, 32'h0, 32'h0, 32'ha300028c, 32'h28c000, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h290530a6, 32'ha414c, 32'ha2000290, 32'h288000, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h24000000, 32'hcac1d483, 32'h1375a6, 32'h31000000, 32'h0, 32'h0, 32'h782f8510, 32'ha61, 32'h0},{32'h100, 32'h0, 32'h5000, 32'h30000000, 32'h5c509859, 32'hc6e14, 32'h2f80007b, 32'h51000000, 32'h2b8, 32'h2f8000, 32'hf4570000, 32'h1},{32'h0, 32'h0, 32'h0, 32'h0, 32'h18000000, 32'hc8d13, 32'h310000c6, 32'h0, 32'hc0000000, 32'h0, 32'hf0000bc0, 32'h1},{32'h0, 32'h0, 32'h0, 32'h0, 32'h8b000000, 32'ha43a8, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h43000000, 32'h4, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h522bc000, 32'h9c000af1, 32'h2},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'hf400000, 32'ha4, 32'h0, 32'h0, 32'h0, 32'h98000a60, 32'h2},{32'hc010000, 32'h0, 32'h18000000, 32'h21d868, 32'h0, 32'hab800, 32'h29c00000, 32'ha5000, 32'ha2000000, 32'h2f8000, 32'h0, 32'h0},{32'h80, 32'h1000000, 32'h0, 32'h0, 32'h0, 32'hc70c0, 32'hc5, 32'h0, 32'hbf000000, 32'h2a4000, 32'h0, 32'h0},{32'h0, 32'h10, 32'h0, 32'h0, 32'h0, 32'h0, 32'h2fc00000, 32'h0, 32'h2bc, 32'h0, 32'h0, 32'h0},{32'h40, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'hc7, 32'h0, 32'hc1000000, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'ha7, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h2fc, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h29800000, 32'h0, 32'haa000000, 32'h0, 32'hae0, 32'h0},{32'h40140, 32'h0, 32'h6000, 32'h70000000, 32'h4c38d851, 32'h142e1c, 32'h294000a5, 32'h0, 32'h0, 32'h0, 32'h9c000000, 32'h2},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h14800000, 32'h298520a6, 32'haa000, 32'haa000000, 32'h5c2b8000, 32'h98000a81, 32'h2},{32'h0, 32'h0, 32'h0, 32'h6c000000, 32'h853af2a5, 32'hbab28, 32'h2905f0a4, 32'h5f0be000, 32'hbe0002b8, 32'h0, 32'h98000ae0, 32'h2},{32'h0, 32'h0, 32'h0, 32'h20000000, 32'h693a9152, 32'he455d, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h20000, 32'hc010, 32'h0, 32'h0, 32'h0, 32'h0, 32'h2ac00000, 32'h0, 32'haf0002ac, 32'h0, 32'ha4000000, 32'h2},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h2a0000, 32'ha0000000, 32'h2},{32'h80000c0, 32'h0, 32'h18000000, 32'h81846c, 32'h0, 32'h0, 32'ha7, 32'hab000, 32'h0, 32'h2bc000, 32'h0, 32'h0},{32'h84000000, 32'h21, 32'h0, 32'h0, 32'h0, 32'h0, 32'h2fc00000, 32'h578bf000, 32'h2fc, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'hc4, 32'h0, 32'h2a8, 32'h2b8000, 32'h0, 32'h0},{32'h0, 32'h6000000, 32'h4014, 32'h70000000, 32'h4c30d8b1, 32'h10362c, 32'h0, 32'h0, 32'h0, 32'h2a4000, 32'ha4000a90, 32'h2},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h2a800000, 32'h570aa000, 32'hae0002a8, 32'h2b8000, 32'ha0000a80, 32'h2},{32'h0, 32'h0, 32'h0, 32'h24000000, 32'h87415482, 32'h188c5458, 32'h2f8000c6, 32'hbe000, 32'hc00002f8, 32'h2a0000, 32'ha0000a80, 32'h2},{32'h0, 32'h0, 32'h0, 32'h24000000, 32'hcb415482, 32'h1063ae, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h20000, 32'h0, 32'h8c, 32'h0, 32'h0, 32'h0, 32'h2bc00000, 32'h0, 32'h0, 32'h0, 32'hb4638c70, 32'h2},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'haa, 32'h0, 32'h0, 32'h0, 32'hb0000000, 32'h2},{32'hc000000, 32'h4000, 32'h18000000, 32'h21d868, 32'h0, 32'h0, 32'h0, 32'hab000, 32'haf0002bc, 32'h0, 32'h0, 32'h0},{32'hc020040, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h2fc000c7, 32'hbf000, 32'hc1000000, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'hb0000, 32'hae000000, 32'h0, 32'h18000000, 32'h3},{32'h40140, 32'h0, 32'h6000, 32'h70000000, 32'h4c48d841, 32'he2e24, 32'h2ac000ab, 32'h0, 32'h0, 32'h0, 32'hb4000000, 32'h2},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h15400000, 32'h2a8570b0, 32'hb0000, 32'hae0002b8, 32'h0, 32'hb0630c60, 32'h2},{32'h0, 32'h0, 32'h0, 32'h20000000, 32'h45391575, 32'h12bd93, 32'h2f8550c6, 32'hbe000, 32'hc0000000, 32'h0, 32'h18560000, 32'h3},{32'h0, 32'h0, 32'h0, 32'h0, 32'h9b4ab400, 32'h15524b90, 32'hbe, 32'hbe000, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h12bd80, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h10000, 32'h3000000, 32'h2000, 32'h0, 32'h0, 32'h0, 32'h2c400000, 32'haf000, 32'h0, 32'h31c000, 32'hcc000000, 32'h2},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'hae000, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h30, 32'h4, 32'h1218860, 32'h0, 32'h0, 32'hb1, 32'h0, 32'h2bc, 32'h0, 32'hc70, 32'h0},{32'h20040, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h2fc000c7, 32'h0, 32'hc1000000, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'hbf, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h10050000, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h2bc00000, 32'haf000, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h18c00000, 32'h2c0570b0, 32'hae000, 32'h0, 32'h318000, 32'hc8000c60, 32'h2},{32'h0, 32'h0, 32'h0, 32'hac000000, 32'h2652a8a4, 32'haadd5, 32'h2f8570be, 32'hae000, 32'hc0000000, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h2b000000, 32'h14aba9, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h6, 32'h1000000, 32'h0, 32'h218000, 32'h0, 32'h16200000, 32'hc7, 32'h0, 32'h0, 32'h31c000, 32'h0, 32'h0},{32'h40, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'hbf, 32'h0, 32'hc1000000, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h4000, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'hcc000000, 32'h2},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h17c00000, 32'hc6, 32'h0, 32'hc0000000, 32'h318000, 32'hc8000000, 32'h2},{32'h0, 32'h0, 32'h0, 32'h0, 32'h8b000000, 32'h174398, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h20000c00, 32'h3},{32'h40, 32'h0, 32'h0, 32'h808140, 32'h0, 32'h0, 32'hc7, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h14000, 32'h4000, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'hc1000000, 32'h0, 32'h24000000, 32'h3},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'hc8, 32'h0, 32'h0, 32'h0, 32'h28640000, 32'h3},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h164a00, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h2c000000, 32'h3},{32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0},{32'h1, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0, 32'h0}};

